��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;������<Ե��a>��ố��PiB���+��� ���Y-bGZ����,MG�gT�����cz���p:@�!���z+bI�G\�Tp����:�o��
I�X�49���$,��N2���̄v���@��'��Ys�PØ�¬�&��)И���)B`�G���f^���o3���k�"^�����=�%F� ź�P�u�v�H���A[T_Q��䳡"�ր�$B�� ���eJP��l����ƾ�)^l�[�|c�����Z(�-H���t�ץr��97�Ǯ]�:��%��������ì�Ux� ���/�=1F�f�>�l}�Jv�yN<�����Rñ��}�\��1�*��+�B�a����3��`a؂z+6R�f%�w�E/c�L�@m��u?N�4�EK"��2H���naA'�.۝���>��51P3̖4���0L���v 0Z��`�o���B�5R���	�/!9���?��D�>oiWi�$�˓&|�B���ڂ��?��Ot,2*��V0�Ճ�Ʈ���\?�U$�(��a`��j��3��h�B�ǝ.�(�$�(<��8��Z�=���N��u���'��sm�X1�}�)#���3#0#�&�9�����pG��ku��%��N�� ���ϝ�('����S���sΗl�P%J���*gcWňx`ܰ(���!�!�v� W���D	#&&!Gh����qV*�>��J/j=Nk�_[��<Q!�h��T��ʓ����M�l��H��ġ�**s|����q����{��@T�yk��[n��d^�2N,���
�.g��u'�}�f�?b��*<-�,� 
�w��/1F� �M�'��gͥ���=�Ƞ8�0dm���߅�jɚ�����������${h*��	m���P�i5��q��U:R*�N�@-I�@��(ʪ�J��0�A�;��b���7�&@PQ����am*��%Erݱ��3�a�!~օ�+�#�p$�o�q�@�xm�7`���g	|݃�����ɇ��*�<��}�xO͏S6�=ݬLd���b�m_xNECbZ�/!�o��8hE8��MGτ��8^fH01�S}*�%K� ��b�$']�.G���D��V㬗�Fu �H=Et����]�H�u��9������Q��v���6�d�����Q'+��>݄���dH��I��yp���h�˵z8=){��|�|������k1-�C?J�Wp����Ox⢪X�Zz*)������MSx�6���/˲�׬}Y�O�2z�`o�j���9����o�V�����׿�l,lȺ�����}��J�ʘM��C��4
�.��5@�SB�O�-I�̽��b�������1���x�J����\��Jڿ�M=�j&E"�~�)��m&|��k'��-w;%�Ľ��N����~U�K����º*��"-к����([?���ն�� ��n�̰�9��;EV,�W���u*aR�U���')�J�Z��"-�Ra"�-�~�U�kA����^r�]Qx��x���\��eݎo��������d�Q}��lg�?�Y�~�@���D0�4C�2��^}���Ǻ�a��A��vg�����GujhBwhT�F��N���Dz�o�Vכn5Q}���E�h"��F"׵��5�q��3�聎ܓ(����9��z���(���w�1*[5�T�4�����SR�
ߛ��ϓ/�]�{V�Ų�D�u�*����n��U�t��x��=�[�i1.W�l"��)l���	=�*H�^v���覸�@Iꡊ���JE&�{3�*c�����VO�M_B 7����/���&�eO�>Gg@~�#2�����D�p�G��y�b`�e�8W�'$. {��I8,�e���En�w=�q��]C~���/o#�٭?��T�@��xF������@�%���C7/��w8ez5�}���y[Ĉ�ې���[%�Xjl`*hc�� 1r�R�)�u~#�-�M����l��w�8u��i�O�����/�����)�����.��Yg��f&��_��x�ӊ#���{	+�x������+TT����tU{0S��cKz�Ӓ^b�2+��Xc�{"~օ8Y���*�:&���>�!�Rડ�&��w{<�u����ksZdZ�Ӫ|��2������B!�)�ûˍ��AʜT�0ϻ�F��Ͻ�7�w8��'�+��Ҭ���0<4@]&﹙�ր�`p`/�J�Ep�}�"M��Z�rp��j? �4���]-%��!�:�X���N%C���0�� �YPk`~6��Q]���]�e���61I�� \�1�lHja���m
�_�97� �N{nL�z6-�����.@ߛ(�.?�y�~�*9ﱮ�3ߪ���^֑  ��8��lњѧq#�G�� ���K���Zup/������B��j%_��1�L<����5��1�����h6��4����O����ל����N�W�gOd����JШ��}�

�Y���s���0~o�͂����z���Ë(ے�V:�΋(gJ�v�4��������5�4�p��@L�OxU�J3���$f_����(��U8���l��IqkDk_'�xD� t<�ES�ɸ  ��l��CAw*|`�G@��y��ϕY,zj�IxV+�q	)n�f��:��V����o.N�ZXCN�7k�d�5S�ڜ��dT�R��
w0Y��V�7O�_�˟��lD{�HJ�;�{���q��t�ls���3#z��u��b���P�O:��t�
x-��qbqj(����ȹmWp�7 FU�!f��9
�lQYvkh� ������,}s���4�NZ��I�öς�~�U\z0(!y:��ə�s�Q�o�X��XAOF�q�ʹ���U|,Ӿ߃�B
8��!T�?W� �q���p �j�Fo�����������DgK�n����|uBT�� %f�Z�th�B��ϭu��n4�Ev��4��P�0��!�o>x��Ҏ��P��Ɣ��.��`�6�}
�P��_z� BmcGO���/kO��k?��9e��0V|��F�q��o+y-#\�Ǜ�(F��x8��������W�w+��F���J����U�Y�	�R��� Ja\���e���|�i��.[��>Ɯ�:;koڕ�ډ�� ;�l+{�5K�6Y
���� l�x�&zҜ9`.�DV�/�f;�A���k�ȸ
�K��U͐�����} n�M��M�B�X�k�����5��I��9�jV�yQ�\'��I�-|�\�&@S1RO,J�C��"qb�X����G����=�5��2��s�}�M+9�ٍ#�[��uծ2@V�Vy1lh��ٸ�4Ҟ��1.,��g�&Vp�LT���\���)G\ʟiJ�����ސ���]���sƆo,�2��+q7�DH�1�Y-n$���@�5�u����#?t���4�u�=r���s$��a�|�}./��h�+�\xι��I^z��h�<x��7Y���^�dCw�Tm�7˻6�$����&�o�tzXܪ'�q-G�*TJ���j涽�y�����.ǜa5��限���o��	p�mp6��d�^�q�3��8�t�a4�t�Q4���
~��W��@�M�	a��?ߢ1|?*H+���	��ۍ�-�H����	""ذ�eF��	��/�߄t/��z������|݃iR|c�.�Xן7l��������bATE�<��cpB�d{��R��� ���u�ݑ�sX9MM*�ۢ�텔4 N4���ʢ:)�zʻ�nl���j�{�@�%�e÷�GUqbzԬ�ۥ�d���v��p9� BW�ա������rUnܸjqF�����#������f�gw�z����qנ��5�K�W�=%�%?�1v)��.��0��^*ʲ7K2�'��ԡ-�� �� ��]��/*7��K���$h�Rʞ��Y�֛q��Ӈ<i`n�{��[D��v�?Gv-�a���i"���(�X	��C��yO ��c��i_�ͤ��%}r^<WHa���V�"�ɻ�<���C���2�]�+d����M2�R I����`l;"���tK��&�+�tlXM9K��a\���k���~/6p��s����b����e#_S��ĺv��Nm�e�*�Q�X��e�3���B|I��C�O�"z�GFT͠������a&)*#q��e��t'�m�'�r�5�
,*���`2mC��lC��J���w	{|F5�$���k)�V����n��<Lv&�}���o�Ò�a#6SFέ�.t�����o��r��ޝ���<��[�8�"@�
tC��,)�Ti�8x"(�'�i.M�mJ�aX�m˯�HX�Z��^���y.`�*�.(���*�v��Z�2�^I�����{Xu���wjy�!����-�q�Ԅ��j���2�j�{�y_��HJo)V�UIy1E9�Py�tk�.���0��#�����Z���=L�ju��9��M=�"�'�F��?��2A�Pcǩ��֒�m���I/I�I����Z{G�d&C�	,nC���&��F��)�(C��[{$�~�d� ח1�"W�}��/3FBA."(k��4IkO�:]`Kk s��{��O�Xp]������4p+y���\�(�$pO�*<K�	�`�W6t
Y�v��}3���]90�%�Cx���f�񦣇W�|f����𩽆u���MY��a�����r,��?���}����O��o��j��)�Ls"��InI�[6����W��#�V���k�Ӌ2�WXK��Ԫ��ݖI����l{ob����7�ͬ
�%�,fٝX;I�ç�;"Ą5�@I���� ���(O^؅���tY�c������4_W��ِ��D�\�ّ�tہ���I��w�-�]=u�'^��ć4:X�;��h�m�l�oFـ���z����Q�	�_�M�2ɹ\0b�#v��Ռ�
W*1��j3�гI��|f���(_�ϛ2�B{�td��2�*�uMm+%��Pr9��a�|e�[}�^�3���Fc�:tG<^��z���>���)�X+�X" �<٬$S���ȵc9,���ݝ��8ܥ��C���ѕ�/H�\���IOq��BT�uY�r�&��a�O�6܊
�:�ܟ�a���@�9�5��L>>�Y]������Ǳraj+��z֠�^�;e�D�D��������#�^�(�.U0nL|�:/�S7��?Ϭd����d����1]����/����o�K ��鐯K��2�3��JΊU�M���룲X�㴡�2R�;��R�Ր�^���6(R]�)�(�A����'�p	��mğ�N�^z���'��Z�G��'q�&:7;)�JJ�R�R��M�;�_���P��g��X�����k�s|��cr)�#���,�V���U!P��=m��yK*n{�:��}28��6��,�lǉ�n��.���P�&ڄ<}�V�_k�B�����E��m�!�a"���1 ���v�Z�>�LPs��	��iE�ۑ��:q�G�BH�3��� _����K��5!tmh-�cFg���6`�ß�)��ȦG� 堤�MQ�b�ʾ��z�����Qo��s��=���4���[�a���@�RD p��hY���$~�P�v���Kn�`>�(��L,Z��l��x}�|���h��Z�s>�q��Z�u��!ֹ�Y���xfS[�}�_��o�';���^%*t��Y��wPCzil2��a�I�n�Ǚ����}��1��w�t� �]>�	j_�� d��Ƥ��V��!��Nw;��^g,��h�"X��`~�M^Y��3{34YN窅G�k�n&;S�}ށf�  ���X���9��X/WZ��z��T��#���[��'�N�4�	@7ݟ���svg����:��C#�G6eǲ���X��)���ȝ��l^��RW��*��)DQ&�������%�#�P��3�6�Y���lN�������R��/�d�zk76bX\�������~%��Є���ĳ븚�ݕ��R�>@�.���v�����U��W��oT�������O��K0��z�S@�!!���;����E�p4B���>���A�:���4�t��.�	CǒR7���2}8&mJ���P{��&�p��IQ�D1"� ���z�ݷgAr��勵tY����I�:��ĨZf�C*��&����n&e����Ddr��J!����u��(�4��6�9����/�@@V�t6��E��ho�-$�ހ�X�k��u����8g�0B��,�Fv4�?�n�rQ2u:Y׭�Q��F�����D|�sbX�N��!�l��@9�����(fS���"�֌���Cpŭ�i/�j$��Qve�Z{u��F,�A8"�IC�����O�yNQ@@@�?MI�3��fkp%��j�����?!hީ������잰�8�g�J�6���:Jս1?����H3�[��3)M6!(�Ր�O��\�0-x�%���?=W�7�͵�V���͞��c��l���XV���p������*��+�(���y"E�1i���I$�4 �#gWEz������k�b��-�����d��-�$3����CͿh`��(�*o��qVk�$pˊ�u��Ќm.U�kdU��x���Ҹ�V*1��Rt�����+��m7�T(M|�X�؝�ol�@�F2r]A��Me����K)&�f/tm��
�����]��i�m�/�9�=)T��M���{A����؁jr�"6��2���+����e(������\�G�6V��d����o
�!P��C�ć�\�ǥ�Փ/��K��hOؘ\]V��Sɢ���|��WQJr#�d(����_Ah��_�i�0��ݱ��ޜ���S����5����X��L�Zv��_����ZLv��j{R$�Y�W6��ҹ���7���&T�/,=���J"�t�K���ڐl�ۿf�/��|��|� �zm�	���>�"�!�w)�"��G�uBh���h)����%���{T�&nK��_�;���{�� �4���f�����#m��p�K �?`Ӡ�A c�0�>�  �_��b9��,��U�Y���{�`�+�C���?�uKXP~�\b��c�ᛢx�\xF��Wv*���s�#:N�GfL�-%�3��ޙ�u>{��_z���*u�Fj2z:1��LS�)����F1]SLʑ+�'�I]�2 F�)��y&<�T�ka�5�F�w���AE�jS�K����{|���P�R�F�:{Ȃ��/`�}������ȷ�f��E%j�?ۂ��mzM��~��\���PM���}�2�S�zX
���UҀ��g0;�j��4y����n�;d}�X�����O�¦߉��+���H�Q"S]m����qi���EH�gM$� � �����.S�8�����q�:̴L3���{B X�Z����WQ��%0݂=obo�D%8����=�}�sA,�����>�
��>j��M��������2��I��OD��wW�G��H=���gę��z� ϑ�Y�����+�1;�[�8�=`�!����Y� r��YMI9��n���Cu/�c�`Y��W�jVk�b���F�sΪuh��x=a%^Q����x�@�QZ�|��w'��Ɂ�E�î閡�wi��B�N,�hK�4=��fo
���K�R`��Z�=��?�`�&��t�k�P�Ǉ��x4���yQ~�w��;�o�,7.�2��,n�JK�c3���s!ʊ��h���E�{��}����C�,�sA��)6ޱ7�wlM��Cj6����*�ɿ�*&ų�9��7��7TM�l�}9����i6FQIs��~B_��^��|j���)����yȡ�%�u"�pb�{���S�� n���
�b�;��QPX��Y�Dbj�Ct�����7��<P����6!�*�&�,��s����?h��J�'l��:�JLI��l��ؼ!���F�!s/ED/d���2�Q*���u�r)�q`�d-�ґH?w?ԅ�=�,o����T��Eg0���
fNhN�أ��>�C��������j�=Ƚ*�h#��L��!x�C� ���=9��n�dopQt��3 "�Bc�t�B*e�-���.D����14g�@���N0��J���v9������Ds,��9�_$)��8�Y�[�����@�����bC�}c���3@s:���C���!��>H��v�{��a����3+�g��a��1�S���<KP�R�K3����-]yr~cP�� �ۨUm��o`֟p�:R��������t��~R�q�7�6��ݭ���*���[<��ɻαp\Pno�Z���B�[2��T�����(9�^��h��܊��A��L����O���|mf]���f�b���1��/_E��ox���~��(}4?�0�0"c)Rc�уC��a�!���X�d�i�mV#a�D�`z0�ـ�Ϲ�Uv���+q��sl)I��j�-w�Vl��z@��Z_d���O&.�^�x��m��> ���9c�~�P�W������cYYD���]i-��{o���7^߁�Okͳ*&b��E��m̞�1���m�[�X�j��
>�SՒN�ƃbJL�+K#���̻�vi�Yb��+���<*i^<M�3vF}G��l�O:& �a@E����<t��&�TaOl��/��M���v������J�K��C�u���;<_��,��+�O�8�J���|�V�=�C��nҫ7I!W4�=�|���.1�N<R H��F�fE��ۘP}��V�y���W%���,�,�{���hRU���|7i��Ĩ�k ;��r�6��'�k5ǖE�?Eg���	н�l�M[�	��u�y��f��t �r�[c������T]a �����ăߤvۋ���Ԫ�UQ�E>�7�y����w��Lځ�BK-m������c��PVWaԬ�a�F� ����o���6ʚi�٧��Tg�D�Z
���q��N�H*ԫ:7�������.��'Iy�!�����U+NC
�buߢ�
��7m��5�$�M���u��i#j����\��]%����}aA�-�hܿe�W
�oUt�DyS��wA�Vӹ�g.�{~Y���rs캗ŋ�h�
�Z�(e��
�0v�,��0��,�����L������<*�s� ��AjY�މa�7������b�˧�_�2k�����#^��ڙԨ`+��4{b,��o�n����l�G7���C:w�ylA`Yk
E�)\��T��o�����li�b�B����N�8x~��8����n<�f���U�h�zvf�+-�EeXQ��jcx�a9��=����G%<gM�����0����l�^`��r���ڜZe���Jn]�OҔHF����k�Ђ��}�fw�b_�	RH��{�����;���������2��Cޒ;��A���}qB�Y9 �.t�pO��>!P�1�o,'��ʬ/���x��.�H�e����%,B��w��޾lx�>�uo��qa��r�#p�c�y�s �Iq���^N"|KI��L�;'��r�3�I��#Ӧ>���h��� k���)����4�B���2� ��ȳ8��<�]7$9���`Gcz�6N�����z�= ��𶩼r.sGL��F�ox��X׼���{;��Ѵ��	UL6o�5o��wG���k�*�4��Û������i���J��d�?�$���,��T�5���o2�H)����"��_a՟���1D��9&��N?A��>¡+`�y�����=�)5<����3�X�C�k�o���;�٢ ���:O6��g�oe�=E�Q��8+���o^E�Fy�R���$6�j�wᣬ���[;�ZS�I7.J�K_�m�Z���0��	7���=s�NY%-($1R'�(����Cݖ����AW�������J=TL6�k�����gi�v6&K��g�+��CXUaw��m{5�) 
�\p�)����>�V*�ޡ^צ�@�$��OI��چ�j� �)JV?%ܜjk�U�#�U��G�RAtgh�ݸ�P�a��P�/ެÃ��@r��i�
9ͤ������nx�u���	���})xÆ|����
�얷��;��n��ú��mN�@3t0Xy���� �}PU��^�{��t�� �����h��0\K��������|%hc���Hk���0�8���PrxS�-��c�m��֘��7��V����v~�\����˛e�T�#�.�ߒ7���з�I��[si�9�MԳ~g=��4+�a���	�H ^p�u�w��w��I�7��/0`p����b�rQ��e��n[,`�;��ܬ���l�aŬ��M!�bl���h��������%����z�d�[m�����C��fC��w��N\�B՟=:��XM�n!Ϫ�mϱ�^�:�~'-Q]�[$�oD����s1�B?��"��f���"�e�ƺ16�����;�O�X
�q|%^JƯu��Lh���μ4~e�h�$kQ�-��{8A�<x$�zg+�(H�W��:W(#N��#�)���	a�[��k��x����ѣ�7߆]�r���S,�����Я�����N_}�x8�_�ֲ�F�R���n���ɄL�Ð�P1����2��e��4ӌ���C��nB���?�0z<�ЁY���0-���s|e��<鑢�����!�kZj���59U�egߘ� 2y8�of1>����X����w�R������3�����E������~a��?4tZ� �Ɓ��9�^x}q��ko�/L�5B&e=�%y=�8�\�Z-
n���Ӗsb��)��c_�K��fD��wbwǈ>V}(�}�r�m4a������=˄\���Y���@^��ZB&�������=U/��ҖVZ6oj#�a�^��oT+�ώʸ�1	hqpk�=`����}�QΉgrbZ�/��dV��um1�ܽU�X�rԺ/�,���"�{�p1�����J��%8G�o�n��\jD
o�Iϛ�j~�P�Ҏ�їp�%�����QCA�I��H&�,,��1�=U�K�ڮ�w�6�(��l�����Gv�2ёX��v�ݰ+�Y�
NS��CtD�QKW��C(`z�yeb�cm���c�c�7&��\�1���n����8d�א�4�TcǠVʜ'�K�|ǌ|�%���7���K�D�C)s�n5�ϒ'��p��B��<Zh;3����{ ��+x��6��R���x�(KP��뒲�q�:^�r�X0^)��#$�U1��Mr�`�.]�i��Of,+��I��x/���#�^�|���>�4��U�p�y��Ѯ�v��_%4a �N	������_��h�w"����ҳ]A�N ��>L���jE�
�;d==FMJФ���o���K�*�����~ӽ�+T�L2&`.���\�+	����<����'^�|x4.�Ֆ��C����t7�k-Ϝ�R���k9�S]������U
p|�A'�;�b�Ti�$� ����%�]e���+���T��y��_���m'��ա�]��(�b�`���*L-�\
�}Y{ߺ�e�
�H��d�D��U~�f���(g�Օ'� ���wꖩ�~W)��h
��Ud����z��s�-�#��1�P�p�8�e_k�s0�r��$�� b�1����a�~��E�6�.{��o�`l �NK�9Z�W8f*j/��׉�y1<�!�QTd���ĒEB��=�>���b�C�^~˦(�$���^[WO�z��r��Ü�>�~�����?���Q]�wiw�'<�n�']�GRYD�.^���>j�|ҷ�#�YT���T����z�yZ��W��`�Ӑ8�2v�î͠��yLC�5Q�mZjB��=VƓ+ߨ ���c-��Kզ���>�@dm!L�����J��'�{����l����<��4��P�u�@ n�d��M>J����f�YC+����4U���M
�7�%�z�Դd�`������'Q�$�C�
���Ǡɾy�1�]nʞI���Yo���q,�Q(T����S ����zG*K���$�Mv����7�����?��x?��e`E:���B��~�k(��:%�d�)���=�������ܺr�H�P^��f�Y=�E�]�В�_>���E�e<��2H�*��ߋ�>S�rg��׌�(0Djr�&�4%H���^"�֌��gE�fPˬ��!Qua���ҵ�gir�ӹ;�G�ݞ�[���{	(����j��V[�@^�߲�o�OY ��u,�T�5���o����N���.6*K����_���C���ĴF�a�	����k�ߐ4	���ݎ�7�UݗN��#�(Dw�bzD]  ��1�2x����3�U�a�k)U��$ەT�eg��rs����I$'<In�%(�ZB!>�U֣�c����+����Ì��!�?V^�a�~DAx��X�I/�A�0r픖��xk����<���azC�q͂e��Rɟݸ9������<���S�OUt.F�R�fi��g2q�[ZY�q�U6�$iT���?v���>��#ɮ����Ĕ�+��6�R�R��1X�54�md���դ�h�'s�R������h�8��Z6c��HJu�M� ���fvnp؜�z��ęP\�T<����c3l��L�>���!�H�P g¤�	����1�l,,TO�R1�������I�3RrPlJ �ɼX¨�0`���v���=�{"4EI2�-���M��>&����@�0�%/i���W'6R,x`k)u� �7]H#�%D$��3�`[�G�O���K&�̆����3��׵���x-�]�#� ��fz��]>�h���D�uV��z ��k��,���4��s����g[ƭ���p%X�J�*��o�|�ϛ���\�^��+�6�v� ����l�0:�t���f�0�,����g!�\��Y�΂��!���5���d�<�@��^�V�ـ�:Y
�|�<�=	"k�F��VR9�?�
�t�]���D�d-�do��z"�K��[�Z�W�L�JS��k	��#�rM����F$���2`9���C["��˗��i}�D��,׻T	t���0��x�6���`�ۍɠ��?ST��`�9Pv-˸A5Yl�%�Tq��	�-I�T=	��&� ��r�wcX���S
������r�
Lݷ� ��յx8H�؀�rp�r��;H),�c:� � �[����=��?!����G���^��y#��r/������?�5K��(�5�����k�r;�E�$��E��F��ԈBv2<D��;O� ~��Y���foG�r�T4QH�Q�ٽSr!؍��c1���]�l��*[&W`�5��l���6W�z涅0�����r�KcB�R����r�I{�U`����A>�����N��)ri��pr�ʢ���\0�y��Au��yw���A2u�8��g����Qܜ�r�@,��H`�V!�hB�e�fμ�Rf�8�p�X�L��?���f�G�6���{��H8s�	�De��Ԋ
5��r_������V-�h"Ѵ�1~�D e^�!�x��@�-�>+�B�����l=i�)6g�����)��(�q+q��j��ŧ���f5/ )�h�� �J���bg|x�,B��.5p
����k��mS߿?�d@rI�-hA��F���|jc���Ť�u�h���
l�/��['���I�I;h��/�?��ݕ��_O�_RK��
-��Q��3P+�f)h�`@�Ǆ6;4�8J��zF�B��g�hE��r{�xom�8qJ�g�3:��/T�}0��l�1��5�a�t~�.�x��Z�̞:���)h��{(ƽw�A�hRM9
�`Y���`h��{���P3*P�	\ak�g2pZ��������}f0P m���Q���j�~�_��p�`nz����B	�E=�<�+͘�~�)������M�-��c��1�� fSC�n=�Z��!h�U��ý���F��">]T�dƊh����Ne^�"dHt�n���o��T��U�۝��3.���P��*�7��G�~��O�5�O�#9Q֠u��ITW&g���3�J�2��OEјcS�,�]L�:����H��75����@Φ㥅И��#�-�z���4�m����D�ҫu��f�rB�o#�xQ���WWp}n)V"�cuU�S����nt\�;�1�*A�/M%x��`JEw_0$MR3V[��%7*S03�
��[C���tu�9��[h��!$�&�4�Q�@�-_:Y����M�ھ���#���.��J�I����x��ewnO!1V�"C�l�7$��1��<���A;�l���U�~���`����=1��"���?�6K7��n�̏W�2�l1)�:פ�ʾ�>-2��R1H_�|��z&߅ɣڜMq!.��U������+�4>�ّ���������:��^��p�'=��U�c��WL|9�7��*Z��eu�tZX~��"�L�,*<��$
0�C�)μ=��8?<�xo)1���5��ޜ���N��r�����r#�T@�@۔Y{�,v�2�-E>�Q=��g��h(�֙�B��wn�F�x�Ҋ�TϤ�]y�X�5�4'����xҤ��B�����62�=�(�����������܈L�óh�̍�֠͆a���s�� �oz����7��Ժ����<ؽ��$M͏R�ݴ[��B��+�]���4!���b0{��	C3����P�䯮e���3ap��C�����1|��C�����
CT���k7iȼʂ8z�m���TWfR�s ���:3�6��HR�) �� -U_�H��]�4�?�h�j�q4��+���_�M1���3���zR����y���|ĂnX:��4�����������	�E�<����Xtl���a���䧃�v{���L����+���ܢߵ$��I�顢���(K<�~���X������q��	�2~�J]9;�IQ�2f75���x����Y�9�6r+����>�ȳ�=:4��0�3&|��C\8�8PQN��b�?�F��P�&0��kk�C����	�>,�t>���B�Ⱦ�&uPx��e��-&W�W��q���[��Q��ݽ��������������+͢�v�f��8��s����}�ᮡ��`UkUd��߅���"��'hݥ�	&�xI��k�`��8kj���r����C���T�[�:0�Aƽ'n���q9�][�:#���L҈9}�N�g6`R���y���pp�gifH�ް�V/�X����W���<��=��
%n�p>��C�/��l-+�X�:vL��ZFtK_��J��ǔ�f>�1x�����hJ���vl�I�� '��3{���ƽ3�QH�0~/�st]f�Ȝ2 R�I
iv���"�%g7��4>c����x�}�E�4��ޥ�;���<�c���sG#�Å�D��Θ�6 %�^���dx�b��p��ሩ�fF%�-�z��t�NE'Ws��6aL��@�৥y�k�װ�AU�B��j�O�d���02�O����z�|ᗒ��R��H��=C�t�}G\���f,@�R�|:Sz�'f��|�����/)Y�5a�����R[q�aʧ����{o���d*7�t�l��)�-�����`L;{<.���&�]|��+�km2׽�[\x��kU���c�"�iF2A����bV�"����Jt7� �"����0��?������+�i����q�H�E�2\��Z����O��p��c1
���>��l���<S#�챀F�g��*Q@��㖓m�)��s����
Y�8ޅd��8��Ov��~۳�H��%�b�D!�h��X�9�N������,�H�l�yݦ@l�,h�P&�{M"���}O�;y���wޔ'wh���������	�ъ/�WO��׳���L½��:�῵}��wp�8Y�*kkp�n�����ӧL!�LUs� ��ĩ�0���n��!n�����oZ*v3�DKtA<��n�5l�#ߜz!-P����?p��5]O-{@AR�����}7T[�j36=~@�:x.A����֣$4�o����������Z=�(J��>^��Z����oP_R�8>���9����?��3l�c��a?Ӡ4$�C&��b9�n�Z�"��e����n�^�=��J3T�a���E0�-.~����jq
�vq��v[�ݦ�֚Aq
�B�P`��|}�k�@N��Mx��b򋟬?�z�.^�ʴ疂
�\����D���n��Z��"L�g����]���2�$�B�UE&����:f4�n��0eޘCjpKuO�k�9����d�_�)щ ��Ch�ɕ���C���y̭L�I�>!�;�Q�_ ���m�XUXiU�zS��1[Z�Z=4�@�bl��`��S7�S�а�l�! S���V��c$��A���X H�O��e���c�G<~���-_����a����Ѭ��F�@DƝ�e��<sj�����ksYZ.���?�ŎUdB�A9��B\�F���r�g!���]���/._fǶN��jU�$M�E����4 8�O�˟��s�x���+��%��V��}����_*�/��y�x���$kMH 2q��{A�wt�`��"��`�@.V♳�t��G�n���ʷ�$�*~�h���"M��j�@�a��H�~��V���FUR��-{*%hۤ)�6C�lk]���F�n w�-�*�x��,/kq��c��Z{�=)��>����^���>�I��:�����d1�✤k�S3�nU���d�[9�8N�	��֮�VVֺC��!��Y$ʨ�JBie��1a�WE����z�$Ћ�T�{�j�;���Xچ� ��u�o�$�W�$+��W$�b��k�P����CLw1���0��^2!yN�(��6�V:i�T��ɛ}�������zx��M�p\���Fv�z�(ӽ�}��R)$c��{�/s�X96mh?((�0�̽S�N(�&�kמ�r48\�@�n��F g��k��X�cߟs��㐸�l$����# ��<2d���Ȓ�~JV���B؜��Tc��*W /�:�$��{��H�B+x/9l�gĆ�Ʊ��T���_H{=@0����]����
(K|�-)������c�T����2��/��?Z�����dL�^�5�f�LW��R�2�5�����ȉ:�,	�py�J+_1�}���Ű��h�؍o�����Q������C���:��ogQ,	7�7q�h'��ˣ�"��c�O����\�j���k��� z9�L=;�e�V�w1��0��b�"��{�%�i6���g7�˪��� �ȋmv��YXx����������$��la�� :��L�����ԕ�V�����TՍ#����u�~�o&�Y���!�h�Ū<-2�c������r۫5\Z�3q��W�B�1�]�����)�@��_�ڰ�����G��m^R��	�n��u���L���x/V��ϥ���H�t�(�ѽ_@��IG\6%=Һ$�n��@�z�N	�$�"�yr�.p���<a�E�H�����bPpE@�V��n����e	b+���`J��Q����1]�ʥ~2�yE�RkW&�y#�#M����5�_﫛����]�����0Yc���39�7�n�a���m��V����%�|.Wq��B/)X|1���k���h��џ~�AC�`?�����0vq�|A��Ċ�q��W8��[?&����EC�3�q�r�/�/��+O�z+������eyZ��h1���	�4��?�y�v�D���#�;8{t�p�G�ŗaRlBi]���盹�.
*$E�4D��jBI���>�3�>�+��mu��\�&>-7��ݽD�8
�I�\|׮j�fEYK����np�6��Ǫ���i=��dY)�� Q��(+	6E��	T��Hq��Y�e�Nb�so�>�CbI����N/� ���8KLV���C$T?/.N��7�vH���(��F�ֵ�Qn��W��jǟ��
�t��Nd�A�[P�p2��U�z0��d�}ҵ��[k�RҔ��2��h\�T��j5�B;{������9ǃU�#�.��#���+�y�����F�ނ�ji�r��o�U�
�VY��x�*6�����^�F �J�bӻp
�3��OӲC�b�$gaF_|㍆q��C�{Zb�*�qLdN��=`���u\�8hkm9��XO�W�BrF���?Є�� "���"V�P:�xUEl�TE
��K[9�>�g,��/�>���rj9H��`N#����銚��A����ʹ���fה�A��Kf�k�����ݭ	��)_�D�ɛ*�ks1m���ኑ����>�*�Я ��]�,�n � �U�J��u�s���Rl��Y]4]0���^��2��c�Q�l��f�J�\\�][����(�J���G�&P�g�N�ʜG v�^r��ýz��'}$�6�g�}Bp���ʡ�M\�U���4ʩ����aO �V������с�x�J�`�Z�n@]�b�"7�Ps��M�'�;�����N�v���Ka�b���Llo;�%Ho� �o8v�>"�jt8`[�8��1N��ى�������K۴,Djf'�`��U������
'��!���F)�����W
fd��w�el���F�Q�l)0��c�z��U��+bǬ� h�nR�?1qу2ؼ��DC"���+�k$|]�9���γQ߂�������N�m�����|tq�z���G�r��?}Rb��2#�M�u�B�+���+d݁cb�<��o��..��ϖg���.�e�ۅ�y]�%���Yu����N#扳d:��9j�6�zZ��y�Հ�$�"Tg����d%��ϐ�Y�����u2��Q�C��7��
��}J;�*N�X�'��:��F��Mw��ʠ��$�3���%�� W�P�1���i���L�;K.����*�nLh�Cf��`��#�Q�Hv���P����$�yɿ	Y˓8E��G0�$o�n�0`A�ܕR�S��,b����J�b�S���D�v"���yg4��$u�	�yW<���j�������HT���f����?A�&�E�$�Al;��
~����E�?���2\C������5���B٤�w!|0Ѳ����-,W9���'g��XK9���9��4�6j�9Ϥ����+gw[��Õbp���5�L��6���=�F×~����!�h�Ai��	�X~���M�P��~0{ܓhG<2��`��e��q�?9:n�Y�����֮��:�On4����)Y����c%1�;���n��ŝR9��*�m�;V�Aj]$�X)�ӆ�=����'��>Sd`�Kӧ���`��6H����O���8�����H���P���1-�Z�u\�z���
�}Ǟ3@��=��!��?����H����4�KoG�NZ��y@4U"�_��_W�-q#���w{�,H���Xv��͚����c�s�褊��Kh�$#�MÄ����ք.���6�=#My�U�Ayǝ�+�\]��)��}�F�P�	c8�����2�^��0��P͉(�?���9Yk΀��Y�;	��eѸg��H2WJ=I_R��S]ӵ�CE2��ӭ���dQ�j�[�`$�]QƘ��n�Nf��Bf�H����`�r)r�)��;�,k������b�p.����I:�h �(�d���_�ַ���0��k��D��������oeXzLuC�d!R�@��ٗ�M'��H�����h+}��c���M4��E*��~Jt�Y:ۍ �N=*��q�ъR*��7��dy�>D���΄�7_5SS@�$�!��r��v�BCJ�.�³�����q������H��-Z�UF�5PT,t���c����H�\��2Sr�Y'��� �Ȩi����*��x��oh�pS��Z4'L����1�L��<V�����~��
�iM�$��N���"��f0ƺ�II�s�̐��MDy�cHk�v�a8,���"1�����	�^���My-�ڹ�om���8!b�>��ul.����<�wъ��=�	� ��uՓ�`mE��ZFG���9�v�G&c����I�a'O�E�+.��}%^����I����=	��m\�,wx�H�	J�R�25�]���;)���Tx�c���V��]���5��y|�n�	}�bE7�� ������>m�խ}{�1��ni{��"�JQ*̲�B��������C��{��jXJ��:�-6Gaͪ�9����*\m38=��������	�\�>T��^�2,����GY��j�r���wfY\��ޞ�!��9��ә��{8z~Q
vǋ����h:X/A���b-�-?}	3lD��z�,��}C2�ctPM�f�+����4�և�4���}�c����G��Rr����׭��Ap�6u�?��uF^{{�O��W�������{�*�l& }<�GO����4�_e<��^$k����cA�[�!랃`0i���W2K1�tE˞!�KI���8(
���Az_<o5���O��o�1����0���wû/�x�E�I��:PpLr�f��\�_&8"j�}"��zk�[�:w0MoDTp�>����!�8��F���
9Ӕ����J31p� ��i�4��fɊ�Q�1D-��p�|Y6U��u��q��n0�nf:�Y��S�PsŐ�X�<� ;B~)���c���^]3�aN��&&v����h��nB���|�w��`v�K�=z�����ub�E��z�L6W�3�i�ej!��F��e