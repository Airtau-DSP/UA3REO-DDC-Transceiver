��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���Ȉ��ݜ�3�\i�ȋV����ݎF�B�0X�'�VÍj}cԱ��e�gŇ�Ep���J����V��p>>�iIJ���R�2���F�����T^��RA��;���id�Hھ�F/V��͞����2T_e�q�ݘ5#k�=^g=�Hfc@�#M��6�@Bc���^�.�}Z\`	wh����<�����1�!�!n{^4@����w~C�� �j�ٗ�3��F2/[�9�n�~L����x!_�����]�1s~O\��☲�����������i���"j+]��2s�&�X�.�K���\���n`�Lb��r���{���c��`�a����ǦR�n�+����=Bone�5f�R�A����> �_u#-�����fxk���1c��;��S?��.�k�p�!I/��w�|�Ō���A�r8��9.R�����hށ�)�\-��>d��������Z#z~��0���)l�����wʒ��[L���P@y x�^�0Rғ`O��S�,���7�i4�1"(�5Yv癰R@0v�Ŀ{��μ�1K`]���)i+�$;�/^�z�_%1��j�f^���܏61M��Ջ��; d(�ŕ�LΑ��r���M
��J��A�����6�k�G)�/|Ƞ�L u�mﶃ���eKC�5��ю��m�1	�{��Ё���=� �U�-�!
�� 5:��/���S�Ri�\^���zDq�L�*���ץ��Ť�>�Y�KK~)ݮαY�oR��{���u>��SX�5��|�\���y ����xŦ�����F�8 k&P�l0�j�+gc|��a�Ѓ��{�BٓI>��FU#u���`�?B6�HK�����8�>���QTΧ;$��~�1��W�3Z���7H�wv|����4�l�x��ↂ����x�1st���M�I����;���}A>�Dk@<ͮRX�յ�����A6b��lQh��s8�ۛ��	Ƌ�k����D���Ԭ�����&�s�#�J�i��.�m�C����y�9��]�Q]��A\D�|-�bU�؜�`�:�v�s�ya}Tda=D<�9c�nE��_�
P��-5T#F��6��c+�NZh�K/2�">�&:�r57�5z���~��D�'�!N��,����f2Ҷ��i�2�|_�=�V峄����{����'v:V�����	Uz�%�3wB>}�O2tD�;6��D�3Ы�β�d{{]�8�S�U0)j�a�V��F�1=J~}�)N�����B�-M\�N�ghm��
d��� b�-�֜�zW�m�k&�+����`�����>�MILE�e���o�Q��|l���������̡�4֛��e�ͱ�2��G!SS#�]L&����!�*��7`�-�Z����c�hc�x3v�`g�����k�G"I�N􈬑�;&n��X�*G��x����r���=��b\D��s䬭�r#u2L���[��vӤQA�#(x��jn��BX#��\H��VL���V�	�D�nH��� ���3s�ϟ��V��N�L�A1�E֖ЊB�
��?��kX���i1�U�/t�G��.&�yv'�Y)�~co5wN��%��lt��e'��s׆��D�q�?��,�Z�/�ZZ�ü��97���_@�t�+�H�!HY�FnN:��${�;Jo�be���K��E���@GA��L^�	��Z-R-�yl̒*�U4,x�y���O%�6y~�@�3�65�И���;�c�'���J�f&�=���t�Xӷ��m,"�Lث�N�h%��H��%���"S�� ��l����H��dEѮ�[R���P,���Zc����kQ�@���1��L�e��اՔm�7a��h����J��Ƨ��J)�4P�p9��Z(��������7���xOD���}�J��ց1e��&�X �sTТ�0gZ��UX�@���?>��^�/J��*���y���R�4[�V�K�p�yw��^�K�U0־�G�'o%|	�O�=s��v����X�xu8vB�����-'���b�����Fcf-�q���o{��^�\�	P�x��F,N��