��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���Ȉ��ݜ�3�\i��4��.��{��Y��?�޻b3;���"�T��b����W�6~?)֙E7K�۠P &��?!f�������\�Γ�PQ';�`J�s�G��W�AA�C]���|�d�I6���oR�_�@g; #ks��NvL������Y���c�[G}�i�a��<i`��Z�	�C? �%��(��[�I�����	n6u[9����+���"����kтX�gZ��.`nm�=��+�,���XL����R|/�%hH�0Q�0�4F۝G�3��Q 	�6;��R���ch���ݲR��$���'��ok����B��x�O�P>t���U��WD�9��C�(|l�7�:xT�^�3܂��9������P�����]�j5�I�O����"IG�ˉV]�x��=��l�:{!�&��rFv[Z��@�ʮ�[�4�P�1 mr��ލki(5��Z�X�ͱ>Iekn=�͑�<^�Y����ݼ��aA�s���M�Q�D�����0@�*�Ϲ=�4z�Z4s�	���C�<ϤC���h�M$����5EA�I~�l�3I�Jy��]��`�'w�!�y/!ǆ���	#�XZu�NO��o*{P��DW�ϮpEp�Ό��e�,O��$�1|�޽>38���`I��?�F4�1���#_#��
���{���T~=�E��=��q��+�hƩ�6�B'��;OJ@��p��b����K�KǯL"R����aC$��g��0�c��;k֝��#kY��>��@���c�U��2	 6�$���?�8�׎a09׉��|����/mv�g���*���&X�EdB���X^�h����+`��c��GI��pK6�9�p��yC��a�x�T���}�� ��k�r���VA��K��Ą}��������iU���\wi��?��nc�Z:).xH�q��1P�k�	�6cśa\'舣�2�P�D�Ec~����>�� ��A2��|U�����b�5���(���{��������z��0|����ì�Ζ���VP���9('L�#)%�\�(�{�����q|լw�H}T��(�OH`��ы,�ú�-�>�u�ԣu�=ĻZ����%�_eΏ%'O+�d����p�*m�x���C.!$�����  F���\AIo��`iX
���@����f0iԼ����%�s�E��!cEc�d��fi2�o�P*����8v�Y��IYx+�C�@�u�s�����_?KN�捱a�2.��.�k���
"Uo,Ig���?�ˮ�"��K}������lDO_�	�J)(��sL̵�m'��6ֵ��EIb�:�+rK��`�u�����ޏ^�$��l!�M}�3{�k��_��C��D}�>C�\%}
Q�#��G>�Tb<˧�N�qS��fצ�A��2��4�+U[��Q��0�@dZ�0ơ;�mJ�e�H��	K�~Ĵ c���>�$�aF�և�߭."���)!
��V'BU���}ӻ�2o�5��~z5`�m��?��t%gS���;*I��2�6`*�<>)�Op#r�:OL�L�� 
�Je0���f,B�m֐��jK+���]��X��9�Vƾ�J�g�I�*=W�P8�@�����맔��z�qF����4n{��=��L��k
����7��t�q��L�]E�'oÏ������[n!q��j׭��9u��ͤMR���� �H�g�d��@%��,�UMtr����НHU��]�n�h�o3�(�m�E����'Y��&�� �+y���h�U��vg*�k���/�3.��%2so�y>�$���oRE�� �m����H����/
<�M��6Qs[_ֈD
57���&��k�v�����	�@[�C�����C��v��O�!�A���>��8��gsPM�	�+{큥�q��3��iU�f��M����@������{��^�Z�=�_w%	���Q�ª >WHJH]��Z�P��7fH�۔L�,m����?:p[�G:�6����>,���