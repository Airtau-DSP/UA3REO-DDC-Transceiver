��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���'�ʞ�~|�A`�U���k�,�ܻ�zc����9z�n#�?Ff��w�Ϯ��^�����[�0�=3i̬�S��
5N���-)�[IN. �b5
��N��@<�"܄Q��X�q�E��?���^�Fǈ��������0�XK�
�7�@�����R�h���������� ����L�!�Ti��hY +��gy���Na#Z�pҡ$���������S����BK�3�W�z2�p����s�[)٠�9ߒ6�� E�16sQv�l�3�J�1={C�:9����ժ�_ooIC�����������~���N
t=O�v�t	��ĭwؔ� ����pʩ���z�v�|z�X~���N\��ZLye�_��t����GQ�R&�潷o��>�j
I�b5en�WyXJ����n�R���9�ЮQl�nW�k4y-}�yV�B>�����i���;� ��DŇ�	4z��N:����j�����e@�X�Ze�Eq�gu�J�*��$�?Fq��h~�A	�ɴٯ{�,��Q%��z�_��Q1�C�v�ߪ��-0O,��6�C^9��O�xiŌ%��=O�%��3mK4�?�ҽ����mgɻ$4�B@�g&��&V��boD������l�k:XK��"��~�� ���>{�S�:��5�f�>�6a `�p(K����i�q4�#�/t��\����@&�JJb`2��(N���YO�H�-J����H��ۇ�!\��+�&��հb���^�p!K�W�x�𹔱�ޝ#S�68�oS���:���N�;mz�*�ov��H؎��-��0+�`� �XSH�yl 3�i�?�e�ЌHr��Iy6
���!�Ql��Z�s��u|�x����
�Cn��U�;�Qy�e23�+z&���o,;�m�.7��Y��o��l�
�8���j
�������o��>�����7��#��w�P�'n`_�Xy�<� ���[��Z�'���U�b䬯3�����i��yU�U�O�m~� �b��c@�T��e�Z�%�#��b�h��>!4.�����Q.rdy�<���Wj'J��*��ۡ�������Z�/�Ҏ#����;!�&��y��L��
���6�s�����1	C�ȗ�L�}�~p,&㵵���GR�����{��s�{/9�[�(<=m��w������Q��U4Xz#j�|��.
��R(u4��\��Q2��G��7�#_�7��n�8T ������u��B�P�W�sq9 R?hϨF[ �?�吝��ıH�@=�,��l�[
*�����r���0����'��%!��a�/�$ơ�kn����H�y�p���뾽�(��"�����h��psF͹��.�u��`�V}	T���<]޼*���AbA��[rO˃�,d�oñN���|�� ����*\*6t�J�YR�;s|˧��l���@A�����Af�!v-�>�o��a
��g�'0u�X/�Ӈ��1���/�����.Y�X����=�#�]6��:5Ĵ�tq�+Y���W�I9C�&{^0ƞ����e$�DZ�_.������ӏ�D�Ң��G�g�%/��q �r[\���o��b	���k?�b��:,H����Ý��U�&��8�|���h��ѻ��#S�@��}@|i�F��.�ݿ/�e%�"������N?�k�:Ӻy�;,O�7֫�3���U�3ڭƭ[ud�bi���¯��j)��"Z*��{�]�ˋg��"�<Wơ^/&܋�`�@3�`}Ϫ�c9�BtU�������O�u�*�G���F��Ȫ�o�}+�m���\OK���/���+�z��E�L?Ȼ`4z�.�@X ���s���tU�R��*|�Dn���S�V�_܀��xc��{�ގ����1��wl�c�^�d���M�C�@�O��L̎��꧴�?6��E��]��Duf�q9	J$��$�H���[�s*����?7�����	�nwJn;��C(�#>�����3=��	Z&�X��N9��f�/nm�$�����A Y,�����#�݇A�ź!��=[x�!#b�C=��X�'���l8%w�DUU��l"�%K{���f>�ˉu�{maݝ�s��͙`0
Ym�5|��#�Y��_����v�J����y��PAE�:��!�����j�WRV0)��}:^X"N���mW�;�A�J5�5��|Q2JBxr�nP�Ab\+��(���[+�u�>t��[A��q�Y�9C�WwQ�"�곆p#o��9hМ���`�F�)�I_Z^ k�i�e��֍W٨t��:E-7�������.0δ�Ykb^��u��>�t8�y5��^��p�Љ��]�2�@p��x]�0o��D[s��w5ajx�N�؅�%�1z�c��u��"�s8�&4�"`����	�̕ݞ���[�b��������o�4�DQI1��Ġ�1��cl���A���lY�*�ߓP���:������z�ӡJ������qF��N����7e����a��G�n� 
%���6zIčm�Y�P0��S�n��8v�$���XR?�݆�V�rO�/�ŞU�U�+V���$H'�����HJ7ls��p���HHs&,��R9^B�d1
�������1�&A5�]\Z1�\^_�TĩQF�a�l(?{9K�?vmRb�X���c��W��<G�{:��4X/����l����i�L���`�Y�iͼ�؞��:���$��g���AR�}L��/����B|ýr�X���e� ]Y4�7f6��Z�)��\�V|����2lv��ҫ�]ǂ/<�/���^�˥c�{Ȫ^�o*h�{��f8>�y	�B��xC�ba �{C[���T�"��Ӷ�
�o'ml�0XɟQQl�V�H�f%�`*��������l�s�l��x�߃��+-;Fc����4�2�(��|~��vgOM~����BH��ϩE_�-��§<���:�T�J|��PY�	UG��Iu����ў�����׳�h-����D���7c�w �`�F��V-3�>B&!��*
��$���V0��n/o�W])�Ǩիʔ�}��)]��s20�I�#��I��0�$�?��®�M�&%,�$��I-Y��a-ܾ���+�J������
^	�kN�G�+��G��Ǫ|R�;����Uft��U3��(a�)�\�_����$��A4��d�	s"�E�G���G�x&s���Y�)����媟�;Ey��ov��2I�s�w�!� .�~�F �v���Z�C��rW�Xr�i����p����645�lV�����yI�`�A��Ӗ��E���P�Z�q�{F��fW}�֊7�qJ�;�=����O:�����S�v�Iܝ�p���;�O�0♧� \>�n�#)�k��$��$HG�ᑅ�s�ve��	��];���Ǒ�4�0�@���f��:N�	 ��;�ꎱ��Ǟ��N��?�Y15���-�����M��BaŁ��t�%B{����i3�cU���X�H�xv��� ���I>�<QnM�g�;rS3/�c@�:^dKt{�CV�ۯ*w�%����:��t����珖N�Å@�42��3���͎)a��Yܿh�5{3ñ�x�����a�e6���j���;JѲ=������~8g7�P.V���?���7GOS���"[|-� �R�n&ńL)fK�"�|mf��x~ȉ��K��u�G�F��i�c�Vq3r�����!���f�֜��Ef�-��#��N����g� U�9��B��N=J1\پ2Z5�eP��Eک�5��X��nW�b3�3r�0�F�H�5�C{(�1��x��hI�:ꓧ�\�3�
����C��Z9X�7Ѕ�ӘH����0�d�?"�o�8Ґ��G�>��/i ���Y�?"�&2�b5�v�j�}"��Z�E��V��5D�Ӕ�On2��q�!�Y �˼)6d �A�����9�8�k�t`�x�7��I��,�]��^���F�2�#���)�,��������O�:F�-˴I4�z�^���n"�Fvq�=rd��O,UǼ��{LW��P�7�W�v_��t����-��R��S'��g~<���n�X~�ݽ�O�7jڳ��m���e�V����
�sT:�M��G�/"z�('�/卣+�.G���p��'˰ՠ���	.g�����\��wm�'�&��F�f���$A��[̀��7��>ܰ�/v�3�w�O���c��ݵ=~ۅ�#>$�yC��s�Yn��Y�;k I���lu���򊶫���ݠd��xjN�俈ft�����Z��cM���p�bA��@�v�a����F��rN�I�oc f*�]�`��:Tcx��Ƣ�ԢJ���:z���p`�T���� �����4D���v�"�nP��C��mA��� +����h�.)v������1	�+�1wi��o$�Hg����w�C3���5���n&��r4��%������E8
�ï)�a�j��A)��[a�c8�s�]kTH�����Y���<3Z�蒦�Z�Q���C�|�Lݽ&�,�RowRï7���t7�IuE�q%����m�.ۅg{���t� �;�oi���ӥ�twK�c��W5�fz��vФ �����)	,����m[�5[�!8Y�?-ڧ��f����3������W�����.g�c-�%d$%�셦��9<k�ߪI�`�/�tP�lFP-%v���=�c�ڡnB��<%ppp~ 6����@���J$M���~1i�q�v���'�P����<���A�<>�9�'�� ���{�	��W�����y$0�~p��=RV���P�?���FXUPe�i���9]1^~�s�_<�'��0�4��#�B�����XAG�9)���|}�o�:+f�W��E�X-vA�w��U�l��O�Zm�AP9X�B st���#��n�[��>C`aa��� ��򆺫������
4��z!qT��HY�TҔ��ܟ�h�o�f}w<���U�>�wS�ݑ3�1���P����S����XM���d�*�!^Q�������4~0r��Շ}ɺIA=B�Q�P�M�ZNz�*��*�5k����u��E8��5�=�;��%U�z���"��3h��*:wsF�*rÞ�;@�?Zʏ���yXD�����A� U�:��V��3vR���
b��B�]�!_�f��LҦ��ܸ�������1���q1������cL��?C��2�ܬ�S�����'�_�d;#���u��S*��3{��Nu�Qt�ï1M�x}�y	����
3��
0���������!�I��N`�TPle�m�W�o�E�f�T)	F�V��t����@jWh�-_ +>A]�,��U��9G��d�%)N�����Z����z�IP���(�
��[{v��E	B}<c?	�6h����U�^�9OF_����Ow�i�8�Ĉf뾇�1qH���@�4��?E�V��g ���?�y웩��b:�$d_�� &n,����=�Ϋ7��n��V���IƇ���f����_��n�p�\c��/�<�[����>n����V'�R��]ȑ��E�����?:9�l̺y�P鹻fy�,�G{č����h��s�Y����5���� ���.gE߷�� vG�8B ���t��gE0k��Ĝ��|S��%~0��h ��Z��15��3�c�\SĨ��Ā���~nk�vk$OΏ`��a��j9X5�����̥�m�{��RXY���W��[ur�����kT���O`]�|,j DkZ̳'L�Q���|؅
rߒ�v8�S�S{��,
/a�����s�ek��f��䯀�?�y���>�E��>k�|�r�U�7K���y�1������Q���s���p�K��"��T�@'��1�	�O6�~��-h���Y����W�6�����^����p��T��0bW����iX8K��D�e��#A�a��+Ԇy�"��
t�����V�N��Q��Ο=�m�GG�̷Z֕����ǄhY��;�Yϧ��i��r+��=o[+�g%��Szqq0zT��t��;�|��A �������ʙu�����ߓ� �#i+��4E�)N��,w���N�I��K���$�Z�G�泚(S��E)�F���o�C��F�����нT=����+����B���B1�h�6�X]�,=��ܭ�~���D׉cļƖ4%�Y�4�7����g�g@r�%�� ��@��NR�(�W�WS������xaVd���2�qm+ǅ\��Bق��q8��'V�l���ٸ�!_�z���ag��K;��
Q��%F:՝ۥd��ɩ=l�9|���	ߝJ��B����ʣ�q.L��F~�G�OJ�8 ���f���lIY�ۓ跆00 f �(��ؚ�����Vm0BJ~�뻛��5����
�fޚ��o,}���a�`�R �̥�e�D�~����t�t���w��k�s��O{�˸*�6H'N��qE�Ȣ������i�T �a�u�̈́���;��_y��^+v=�iW�0����BV��Q���I�!��+Mq;	r	�� ����_���������2�wȄ�)�P��'��,��X�K}��1d91$���{-%}y��_���1��T�Xs��W�"��x��]��k�e��VS�2ud�6�t�b�a6�c3lr��7��@�?�� Jr	��BB�!!B9Y��W����S�	O�X\@I=86��!��dU[a�R���