��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����ս�Mm#�&G��BaUG����5R�ۖ��Xyc��N��2Wv5�n�[��|å�6糕�=d�����Q+��4��JiVE4I"6ya�@�Fwɮ�V�Nhݽ���5Oߍce#�)�<o�]��ͬ���T���P���W7�}��{������[����qG�*9C��~٧���ͮ��|O��:��)~ �ʽ2�+�Wȿ��� ��;/C�����K�}QQ-�8
H:�^�p�
�s+̼F���2�9���}lb|���|��$�\lq��q�ɽ)�6���1;2���kG~z(��OGq���R d��ҍ�e�5$2��?��#b\����eT`���_.��o�1�Q�q��$����G+��E<%���7C~w��I����K����X�����&/�[f��.���ڬ���stܸ�1}rȌf|��0�����/�2�+������ĵ:�{5/�˿b��N���ˤijgҙD�NK8�?Ue٦{�?{>�y�S�E��<�0b�2��8J�'��gE����/�6�������i�\���N�wh�i�=��5Vb��ύt�p�:5so�Q<tM�i�֔�E7Q�J2u����	x�W6ҽ��ۋ@�6����t����Ta����ٛ�����w�簗97�L]`_oP��5<�|*5���\"X6FWD|.�m���)<či�d���X$�}ӫ�����mԆ�";^�A��]s�tT�~}�����N���Y=cQ�p������ݽ^AA���6jh|�;
�b*�B
���ﴘ�+�Yo�ɈB�/�@�{���|��@Dʗ=�����t�Wz���4Veo��g:�����M�_��ERA�DaU��nS�)[vzV|�:l�/��n���_�1c	
��Isfz�{�61�cWDC�{f���y�<'D�0�u�b\�� a���2Ϟ���<�5i/�ܹ�>�����?�μ�Jc/�Y�tW�������ʔ���C���Y�4��|qd���c��/×�o5��G�>�����7̘��h�O����C�x_����ԸkG�F�ͮ�'򸳿e��£�B��8_\����$��+d�j�8::a�t��8�N�%
`��mX�� >�2-�^=:V-Hh�#����9��v������.>Q��c�g���t��Y���D��a}T'k��ɺ��f�Q\� n8t�`������_<V��u\�6����-��C��,n���;;�Բ�x�2xQ�OoW��1�7c|/	[��y\���S��1�g)�i>j\�U3y1L	��#%���K�29�OdK���5z�>h��֨u0Zt�ޓ9�(ĉR�l��eCx2G�B+�[sC��HEL�����vKR��e�L0l���B�/���&�b���^D�Gk�����A]��of�<�k4[��^L0�B�D����6�����~����$5�P3���8�QD���2�9YS��hzh͡#��J�kh�UCqyq���H?���O�M *�H���{�@l�va[iL��s��R��n�ӡp�˅�
�`j7����R�N}�:-e$�`K>\mw�^�i"��y�?"G�$70����4��0>�>P�-"��Y�lh�?sܭ%=�D���Ɲ��[d��������%f10ߪO"/?�P�岉>Dg�~�)��sq%S�Ӑ�q�!��ehL�K���k����EX��������g�S`ѧ2(������49���b�2WP��v����cQ.���$�j-�,;u76�(�ӫ���e�|~�5��W��`F��I�F���mrs��}����c�iͽ���a?B"q�H����,�[K�{ZO�v{���E:����(�_&
SB�7����Y5<�zl��^��n�W�����Bh�,|���)YH����-]�hQg��)TG�(���5�ru�ߦ,+��v�=�(4I�� �U�d>�%�M�
�������q=�Z0<=l0�� W$�<���
8�SJW����3�5��H��]H��`A9 ���A� 7�6}B��FY�΅����y��x9�*FhLX�V���n�\�:J����0�htd4��4�ZQ�� R#̔�؈uV�M�Y�Rs�ۍ�����l������7�\�T&o�]��vǜ��2�:�ʦ����0 \��`PWs��7k{�x?����7b߈�y��+(�Y#��	D��"�[o�U�er�Щ����iSȂï��pG�h�,����U��9D�ջ�[�-sT{�(E���q)bcB�r��_q�F��ŕI^d$������r�sF�ju.E �o�V+��\��k���p�s!D���/b�n!���=G�*<������:�^ J�\|�v�=���3��f�?�$f�'���3����<�
8��e��9��=�
]�>�c݈x �����@��f���C;�D+X(���e:4	�L�,����S��YW�s"!G����������iR�\Ik�/��E�,g{Ĩz�.�&3�[T39Q}$�f��5���� �G��Mr�._(w������ _~��y��2����a�ݼ�!�-�`����.NO��S璂���6���G�ڧ�w��xCiT���l>Q�n�|�ӴVq��	��u�}S��|-�Wݞ�j(�>h�?�7�S!@�3J.�~��&���`6ڇF╌���]�U�u�/6CAn-b_8�*�-]�<.FB�!��	�!�Nz���TW(f����,������'Uj
�����.œ-���g�N z�W�M�m�7$�Uw��,}���(D;���toă?�����(��3�N�2�C�� �`3�'�Nf���s�^��^���ٯ���P`�cg��y�b'p�A��EQޫ`���e|�8���{J$��ߏv�א�]�h��&1��&��"�����$
�/�5����P�A�yp��db�ȷ8��T��&9K�Ha�^�4d�94"�86��۰��u�(I��RfټU�گ����&��G�8�R����\��=]"�0*���($X�4�r�)�'<���8�L���D��!� =Ksz�)�|�!�oYH �-��G&Q��Û�H���r�Z�=��q�������6��{gَ�ѡN��E�P&K����ٔLU�����E	�]���;�|�WEi�������Fp
�@��+�/�Jb+4�1l�t�
Sjĵ����Pn�����L�vM$ѯ@p���|��0�Z�栘&��$���^c�o͇�l�$�S������Ȇ�߉68�LV����YKP�J��<���jEk7K0Ev�G2.�_��x��jk���PaY�>���j	#�+ә���5��/�9�@���G}�Ԋ���"�֧X֦�0ֹQ�tX>�����= w����I"0�z}�H�yڔ�c����6�|.6��n9x�� �T| �Y�����O�-��$�Z�'������e1r����Zn�}v�M'ԩ�5 =�3����4�@U����E�n��w���Tե�[l��̅Q��̽Cm栘��d>d|�m�e��8�=�{�|Ű8x݀B�yT<�Z8���[J��� ��1N�lQOL��\�k^B{�h�D��;tUsi�P��.C�W �:+��1}��}g�E� 0���i<�:3y�>5�C��4���Sʏl�	����@�`?�d�Pxa䰙�,
�>4�
�]�Zof�����f�Սb���w?ָ���H"�Aj��ձ����8QW=�y�/��L��������(���j���նԵ�ܳxdGC~( :dpqcr��#���}��ET7 �k���'Z�'+������xq�s,��CLݡϊ��b��oU<�@60�q���F�Ul[��H�<Aq�Lʐ�\�JM9}�U���PAX3N�^�;�����ɳ� �1j.��YQ�H	��~V���T|Iz�%c�����՚͂!��o��������J�K�Z} ��~1ٶx�F����YLs���׉��_�V�e[ʧ7b���TB�2�!������]�����8ƺ����*b3k�v�m(h-	�����|��0���_nz��:�bY�8�@8F!�����7ܫW�BW��ߚxC��� ��9��b�`eY��&�'d�U�ǽ�J�
Oʔnm��z�@;as��;��(1��J�O%g�0���cW���a�KD1��-��<����sX���CI��3�W�����+4�n}[�?�~�;��	#�I`@��L��q!�B4�,��\T/�e90�����P���n��[-�r��n����UO�&�~�Ȁ*�>���w�9��bK|�4�yk���SQ�����tި�M-8�6��݋��&Dgm�������:JI�ާݞZF��7�%�d��w��2�H,�>�O��*����Ho��M�-� 1d�3^h�z�^ S���Gysp�<����+$[� �;�s�^��(�@��[Y�H/<gԽ5���9,v��yKi����w��p����_�G�1�s��M~�K���B�8"�C�8�uU}x��8sCMy�<6����	<A���R�'���v,$|�9T\k��KP��@�Ո?`��*^�Gï��g#:����=��-܅��P�6�4:� *�� ������i��^V��lv�D�ƭ�Z��H�X��T3�@$�_j��o��6_��l*�)9��N�K�{��&c����O8�4�p�%
��/�!t��������{�f�S�B�uz���p�z�鎢��y��JD�l��ִ<����UΛ�$z���K��4�/٠�V\�]xzT�g.Es�v;�T���꞉��N�n�>�PQ�q��?w����-'-h�B��~�B�j_O����W��֖���phs6X��v���������E}eԛ%��L�K�{tڥ��K�-�z��\7)�F:��z��g���?���ϻc��a��Uz�A�����w�V��)��5�*e%�݁�tn����#s�4�^�m�6mG��5sM�~/S������4�� �ţ���@�����a�����lH5���H\���֑��"�J���Xu'N�e@��Ϻs�|�}^l^�ZK�����ss��g!��
mD�@���'4X[��X����&K��[!��l��ȼFM�E+��uˏ�����"O���f:��a�Apk�ZQ��p�1=�.����AGۋ�EK[��\����4��f����=/�j�� ;ۼ�Hհ�@��~ΐ[�A���R�F'�^Kc�Ǖu�W8F��G���b�U�~ ���h8�~	��U4���B���Ж֩�{�,�{�������ubHz?.�,��>R��o�V��Զ��.ޓ�.|��>��̥��M�y����7L]���y;���W^�\H!�|��T����\aL�fD��2���zXx�b ��6�^S�r�e�&�Rf�Bs���������~2���"�����C\��ۚLYo�V�:�q�WT���u|\w�6�f���u��/O�^¦;\������U@ ��(�.���p�8L�ÆYH �����u@��e�S:笉�\t	Yͷ�^�evJG�/�շ_&�
Oӧ퉕�ڕN�WU	�g,�n\ѡ��JK��O�B�o��- :K�Ü�㋿o_� ����I��^�&!y�,giz���Qt��Ao-y��"o`w�	Mc������M��u��"G�7�1&�|DD����w��
YF�"�ԁ�T����,8�]�Q6�����ƫ��G�M*������\����v�Nn[�9�\��`s1>����zVk������EHH�Y��7���V��y*��;)U��A���0#c��~�Ó/F����u�@�����\z���uL&��yۯ��X
XI]U����߹R8���{2�s�Z�ob�,����v):�g�pqVaW+2�=l���}}����ӇƵZb�K��d؇���W�T��:l�qv��W��`��I��ŧp�-$m��Z'�j8)W��Y\EU������ʌ!y��"�Hf %���-�O9�Iz�����؛ ĊkDU�=΍y>`�ZaW�z�U�v�]�]`�� '�������nW���A=T߾fZ!��n�,"g�t_ߚM�]�br݊^�a��|,c���)���灐��,�f+Q�=Dp�@�Y�޴����p�}B'ܸ�b�%�谗i���w���r�ʁ���-t,�nD4V�yĈ"�����3*���L	ɥp=�5Q���r�@��Ҙ�OJR��N4(I�� IO\o�t?-Z��\ ��X�DHgk���R�&��c�=���ا=�~.�*���.X�W���)��P�5q��L[�a	�����= �x���Կ��U��p��󛿳p{�P�z�I����v���i�tTH!e�
Wda/)|��ē�1<XCM��#�=:^Dlι	,�0pES4_�4n���(���nv�� ��g�dfm�ة��A�yƒ̯�-�l����i�m���c�wy�ؼ�ñD��H�+5�r��!qg�]>}��EQ�vh�J	�b~T�RVad �L�cԮj7�E[Q��{ڰ��U[(iǋ}�`H<�*�q�x'v�����uKa��K��ܷQ6�bdncO�SOy���/����Y���&��@j����:���#h[��Jr�3�{��*J+��>��\1���Yڟ\Q����B:�P�sg�S�c�絡0&B؉�S�G�	�7�mU���'�.Ž�,V�f��V~����`b�Ļǌ%<л�rD��3a������e)ؒyQP�`�mK��d�f��Qjd��8_jN��8���wK{z�<)�AδS�	�߶&�� ���E(�s�usrL�~ո���7�'@#��>#_&D� ����5 q���!�����Ruz�K��)in}�:ч��\-�Z%�*���hiv������HW*C.��f��9V��Ot�jU�7H���Ul�Aj0b�:�&�{���+x=��l�_SZV1��_��� �����YThU���i�y� 	V���j�&!�	��z�饒��JӾ�P��5�f�w�!C��O*��]-^{����l�Q].�$��R��5=Y�'J-�Iѻ׆���|#����!��rp@�9c�&I���8RK%������'�Mpƥr�k���2��i]wr�Gj����jvB��{^��F������4���X���i���dEj���O���4�����h� ��Yp��t��E����Ƞ��NK��Ȯ���5:�|
:�ਂ,=��P+��Y
��U�L[��^�5!:𹏤�������4Lk;��6WdQ'��C�R���<��>+���C��n�"ϗS֫�4�.��r #�{�q�Kwc,|�=6h�	�>'̠�)�(�0��������^ꮇ� 5��1ܪAXv�9�ay�X��r�*+Hs.��\>k�����2�9�W�A����H�q�<K�����`-�n��
{�u#��^5����z����u$�U���5�e]�|Q�r�����c���wo�c	rĖ���ǅ�D�'��`��c+D��(G����84��w�P4ʹ'Zkءt���O�k�\ƐjvDA�z/��.��if
�����k����va�V��v1��S���i�����e�.���a*��'S�L�*bj��ڄ���*ĺٞ|@"���Mb�b�%���K�GGp�C8�Z)�J���l`3Ώn����&�&v�k<��놕�(/�6Ap#&u�Oˎ:���4�ki����֯Q�.u�C�Q��}B�M+k�(��Qi�1���	Q��?�LB