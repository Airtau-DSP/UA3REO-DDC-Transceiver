��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k*(\&��Y���z��;����1~;ó�!E7+ Uߟ �v��M�a�v���]�P9�Hq��;��p3��W�Op8>��N՟�8��i�yM�O6
m���h�V����_q�
ɏRa�H�g}�63t���&�X�~�^cȮ>�!����;R㿆�UHd�D8���5���_%� wt��fD��z��E?]Ck+������?�]�O�q�W��Z������B4]��m\��?�!�!�,Fv�����$�Ti���]��=k.��������CE��"ߗcRۢ<��!bn��&��.�s��H�'��:��v��v"��M�ŋ���zl�[��� � n%X�e0���P��Nz��b�H���K��TsAO�����M񅔞�R"UD���ͅx�&+y�I����F���A��.��$#�}�	
5l����Z�Y5��|��X�gN��^u��2W��\�/�c�i�bߓl���F'�IC��nRZ�k/o�f�VD��sJp��J�Y��q*���xFB4��#�%���]�`XZ��ɧ���r�3�8�����_�R��$'�Q�Y��F|`�+WƼ��L�劫���?��}w��Ϲ$��j/�F�D0�g
�ͭ�t������M�O��*LZI5:R�+-�����F��nL�Җ�f�rD�B�sV@7������O�������Q}�@K���#J{�@���P�d�!ϱ=�ڑ8e�V�w���F��Ad�u��Df8dZM�t�Ϝ�<-���J�uOVH�B�'K�/�R������s��l�ifa���#�d!�&���BA5"�����C|{��߫��6������A��>+�cW&��|H)-2`c����80�nO�c�!bQ�o0�	mk����Ɋ�AV���(w�N'�r3)-�P��Q���|�sg)�gJ���)�Rjۈȏ2�Al"���x����Wu�(Aq�?���1L������π�\���z�zꅄ�	?_�j��Br"���� #�D�k����h���)�{�g��@�zB`�}�lZ%￀m�Z�Sp�~@��E����1����r��AT.�rwѥ�T�_y��%:��$�,�>��`�D����m��I�Ĩ��[p�n��b�?y�����#23F���:D&iT�GU�i�t\�-N���<HS#80��_@I��5@F���.� ����F���<������*�%���nI� ,K�L�b%�F��#>�Qֺ��i6�0��L��C.}f�E����S�fn�������?|��>}n�9N�o�׌���Dܲ��d�p��KGJ����5���a�� R2�a�pq�S�M����N��
�������>������0'�' �;��ھX9F���%6�XP�����Uvx�IE�ҴT�n����	�%C�G����o(`��w�o?Ѡ�xtW���E�ֿ羽�};D��h�6����� �����X�QAU�ׅp8�� :�Z0�7���
r]�����n�"�?^��Q�I* �L�, �-����.�����TH�5��&{v`9�������)1��j����&]Poh���Q���K���2�e�i� P�U�-�.����]��k�{o��=�n0�����V�DLp`�I��������fV����q����0^���!aŉ�(P�D7�`��t���,����讫��>B�^?4��]Q��q�JGΖ_�f�ŧi��d����v�eސψ��V�~�HL�u9h��jvz�O�����k(��i�w�����+Ro˥��?%H�D�W��]=��%��[M5D7�>	m��_�����r�x��9��w_���\X4������0^��.��u����r*�^���=F-�<��O$��D�����$��=�h�BD�q�@��hU���@�<�JG�Pp��n�̗��[8����ΎwVNNz�g�������m���dk4��^Kl]�R�_��F��qx��),vc�)�3� �5�"S�2o�t�Q� ������]h?#�W�� I��Vud��Ä*�2<�Q9�v捆�^�W�O#�����{��nm���C����e�k[c@�3�=*c\���{�(�xY�+������~�g��(�\�ق~���\u$�o%>��dn�l܊,�a1��_�7�'U�檔���� b9r�42�/�?��m�CH�ʹj�`X���c�+��o!r@��h<"�>B-�	�Ed�{4�]l�ޟ2,U:	�{h9*q֨��Ag�}�Q�`-A>Wj��������Y���"n4�O��d���,>W!�R���5c���]����߆;����*��/w�ϟ�{0�=�O�n����7)U�嬶���F.�K=�:�p����.i����Hۥ>/��GL����R �Wޅ9t��D
������X���|���_�,�䍐�g�'��Ggo����pKm��w����ޣ��,uQL`���*�Q��H2-�#�v��)
�"%m~v�ګ�2)U�愠	=;�����o�CƗQF'��Ӯ&�KbГ ��B��sa3E�t/�	^�e�2�[ȩ��Qb��!W`\%7�_%��S�c��ñ<��l��'aL� c�����˼t]=|������e�ڳ���AlWfc� ��qe����x�h����i�ܱ������ r�x�oh
VL1L����<XnO���i9�0-�F��$���V�O�N��*@�&W8�ϩg�����e��SQ�\���hMͥS^������C[��ꪤG/��K\j%����Ƅ<A���̹i	�����<� D��{��߃Er�I�����}X�գD�{�y��۴-�;��۶�g	���9�i�m���8���u�;��y�P}�p,�]d-�g5�o� ������.��,�Kx�#�(/���*)���[��7��Xwth��n<V�=^���aX@mP�cD�e�+X�a��/&�z�n6d�0��1z'�)��'���݋�L���15 6��޳� v��hɳI_���A��a,�u/�ڦ�*j<���e@�&U/��䘆{��X.����r���/�
�'D_�͞?�k�P0���������t��<u��{v1�W}yZ
�������� `��,�������l��[q{	 y�;��ݞ3r_�F�V�f6�#C�<�"��_���`@������b�j��>r�?�sî4��&Xl�8QS�p���P��������.��'/���|�i-��D6N�g4(.�O^��褾d<�����Iǽq'_���z*��6�����|z3a1�ӌ�M����Rk˹�#zo���"$>����M5�HA{�J���l�Ż+v|�8��=B�whia8�� G��[�s��͐��3�[�D�z�ɬ�����6��ۇ�{�I0�S���1�Dk �&V�[�<�Ā���"�����z�j��uY���(��m����]���>���Fѐ=��� :�0x�e�q�#:�bD����;�A��R�#9f�Ϲ�Z�c�����;Ͻ���Z|�`o[O~Dy��j�ʪ�!�t-�t��nE4�*y��L�s �d��~��y�A.�:?S�a���Ʉ~:{�֘��20�h=D,'�3#��Q|5R߯R[\�F��W�m����&ݘ9w'.��R�{H^�$�;���e��Q����C)��C2����[ƪoo�#������L�Ҵ����d����ލ�b��CXvi���/]�S��,�j����h������ҫ�f�ns��Gep�V$N��=�@���X��+����kQ��	�_��p��w=R��g��4-@����e�/��,g��!�D����_�V%u�1!����vo��c�����O�!/���8�K�Y$�C�ur+Ti����1v�k���G�THU���%��˿�7���П����c���g��["}��X�r}��������|�\�w�4s:��="���"��1�^}��� ��)�]:)�F��R7���G�Ǡ����D��t���Vw֒U�b<���Xߕ�#��o���\B$L���$po�`3E�$c��5��x��^o��=Q�bΉI �˘@��������Ҙ�,�����}�\˴zAN*��R��!�WSu�Y��she(&�]1�"2�'��x�R��C1\G�J�U"�<R��Cʾ�7���ͽ��7��W"[CE��+�ܳKQw����+�S:<����4{�=+���A�ξn�!���T��,����&xj7ۛ��=D��OW:�^{�p��ǡ�넲&zc�8)���ڳ�FI�O�4U0���<P�����,�4�
����e��͑#-��\?�k!��+8�~^�`w�$Eԥ�E+6:nY�&�I��ၥ��ٝ��E1�1�d,iD�����qF�N�(����cŐ���*la1[���8�l�/�7a�(���F3��J���d��������l�J�`cRh��5��ee,*���~O�8�&[�� eo�>x��'�m�Ȝ�#���B��bH�Ϙ�D���}���5jz-�'(�}�c;
��]�'g��<c�����Wj��,O���a�A�T�9^�Sm�*������X�+%�e��?�U�(��Ͽ��=�p���g�]�a���'��X̼��%w{��W �?�N���>��wQo(��z�M%�����d@���X{+���i\f�Rd"��t�ͯ��o{���VA����?��ap�Y��Q[��i�	�0Qz+�h,�*54�������7T��N���KV��]�����`��<l뚁r���x�����I2�ֽQ}zU�6fW��p���<\�_���c���/���7�����z�����s��wE#E�5�{`�8�-�ێ3�Ǐ�>&&y�y��������D�N{�ؽ�]�H7�c$Q./9hJ�8�k2-�m��~[3+�y0��"AЏ:��<մ�0/�4zy��	��u��s;Gy��j�e���p߈!�$�x����=Bxx��yT��*�������u]�巟��*,.m�d�ku�tc�;�`
���#}��n�*f�]��XeT+�P@U?X36��;J|�`PJ �:uТi$H8j���n�rJ�|�%]7;DX��wAN��ȎAFJ�q�n��K]M3d�D%��jUx(\8Q�Q��KP��0�x�����z.V�`�N1�q��"�W��	�w'Yj�a�t�i�W�Ƣ��R T3D��s-.ŷ�
��vY,�M�ys��3�Hs�1��c
��kJ7}0�>d�I
�=ܒ���Ð���ZN����L��~

�{��v��L�ᙡp݌���_G,�-̿�l'�]�5q��p��'�|��o�j��W�s��S�W� ���(�+�U���Oۼ+��'��8� Z��6IKT^��3����Vd95k�e����<;Y喲��{�݊�zc�/j��׶+�Fo�~�{\MK��'��j2Z���3��et^�uRQ���X�NK*8`Xn�U[f�kpN�	FVc㥈o@1���4�#��D23�^���_k"��y�ZD�q0�%��2Mk:���fE�]\y3�>�X�-���.���
���EF�#L��JVQb�S}�_���^�u�hnބ'���K���xlC����!\_lٟi��%��۞U�Ю��K��F��T�J�q�\썐�%t�j��}��7�N�+��Q��9�UU��페��s@Ōp{,�!���w��EF`��``B�k�)�
7Y�M��7o���g���B�gvv|��3�e�����s�=�"�8�����$!o�˽+�j���ޘ�R����́�����������LM|R���ɫ�V~Ԧ�����En8
	#�)����)d�0k���3&�]��}�[��%��f��Qe�C�YD����9�7w�{����Q���Ei@8��0�-�N��x��_�=Ti^)EU˃���OgL�'Z�����>�7�3�Oɰ%�R���M�,��L�O~��W��(C��p㡻]	ט�>-�I�C�����89���ߒ3���O��H��0�B4B|=����
d)vq�M{�:�l�����%p�M+��*r'j��%���!UE~.��e]d�;֭٬ �BU!S���p�}^���xVqL�W�����Z�£���x���(��l;��Ċ�ϛ��un�U�ñ������K�&���
)�*����؇��&Q��Q#سg@�6%�]�#����y�����;g� SL{a\�f�����+O? �E՗y9�4K?r�́HMv7%f���MN��">H�v�bZA��A����h�+`��x�p��8�f��j��(��)�7�c�>�!7C�3��O_�����s�K���a��Qx�~܆Უ������\}�׺D5�N�e���)���峃��(3�E������K(.r�u��(Q��	�UT2SO���lUPZ�2o�����%��9�U>�� @���m��Y*�^��f#�5�!�Ţ�kkF;oYE�=��}�3g�~�0<�g��K������o�G<�H>���r���.�^�9�B����ْed���.��yMC`�-t�i�3�����zS?9$<���N;����i2��Z!�d������x}4�֢mb+���E�S�nxw��u��M |�9��2�A,���̩vK��M��+\��� ��G͐|����	�ae��]������1�z��7:"�~Q�:��*��V-�˥w��}�F=�|�����qMo���r��Z������u:��ZE���܁�X��#$�`��8	�6I�}5&� ?�i,�6#�V�8���d�4�}G��4��^��ܜ�����b���"CG������F?���=�F:)?� �7��y��R�����Fr�|�C�N�>.�L�"�F����e�}��@���L����!���.�����>��4���R�E-GF��M{���z�� ���Y��m@>X�"���4��(�Lg���j=8�ټ�f5O�L��?�t/K���#70���0�t$Nk�=��fjfz4x�+�����!�b1��vl7�����0��R�U�HRm���$�7I�'����E�4�F.X}��p�B���V�2jRA�,�V@���z��6aHG0D#f'��ɦ�P��f��&� ���-Q��4O=�3q%��|�k7��k̒F=ɴ����*�c^. vc�v��sv�;64���oq��W���=J����wQ���,��h�eٜ��FtJ�}A���M�M֮�
Z-�y�VN9bX��j�ڛQ�#���HJ�\���57툎���� ���'�;���3��Ev�X��|�D~�����:�]�\65�	|nd���uv��