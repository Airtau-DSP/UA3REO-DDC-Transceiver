��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J��%c����~pIbX�˘�u��$.�H�F�!�'���/����|��{۴�=�\�����qT��M�V%�킹zC�h��P�R�U�#�sR>��*�GHNW1��_�Pό�l���:^V5_)|rg�%A��j��<oH��7��ҭZ��F@���s�23�o;U�����'�tȬu=䠓�mV!�$*�Z�oL)���/�s�?���;���&A$�K�|%�k�6�A4��?�I{��fo,�zEC#�5�61$��>�$�!]�.~M?L���'c��z�񜪤e��J\�>S�SZ�.��u9�'����ҋ�t\�Rt,Ἲ�>��Q;FF�LF�j�:����k��W��y�e
�!�4�܋�8��?�-Ԕ7� ��CytrZJ����
/��C��~z˸��ٷ�q�:,l1��KJ �I茕Ji����3�G���l��S���T �����䍺6���.d�6�!�6�$H͇������8<��svū��A%,#}#Q�!<Ԯ�:�O,؇k���A�����C�1O�Z�(�G�I��f�Ћ��^�w�Ph���b�s|/{>|��m���3>���-�?���#���S8&H��i/0�z��.W ��9��v��m��)��n g�@$i��de��a̹0�FCX0Ů��in�TQȦ
�(2K3H�QD�oǬ��<,��p���\��_�Pp%+vi2���O�o�M���QI��K|��5"����d-R�9�23^U��S"U}�o�E� 6,TXy�܍FٷՋ�0�l ܕCf?M$��Or�˙�'tO���TO����ˢ�߬og�K>�j�9����M�jdX�g��s����d�`��Q���|IhIh�	��ؿ����oy��� ��`�,:>v�8������O3�0�G4��'�	�z�R�4��K�,Ѩ��C��s9v��Q��Y�vI	o�a�Fϒ2����6��G�9j(���>@X/,X��UB?`����77Q=S��"<�4�0��$�;��
����`�.��j��!J�ݏEڐ�דJQQ�[6�a��^�ij
��`�<^߾�aUؠ�������4;���\�>�l�7�} 4�2rl��5���Mŉ$���1�Nq!v��0�{\�n��~D?B>�aw���CY�xp4�jx�¿��I�K�Mp�4�ɢF{\�nQ��i���d�E ��U//� �)����v�Nk�)շղw��I\�W���*�F�� ����)����ITj�0SD�m�Эܲ0���G!���("ڑ��o���J
T�q{����/�x���%v���Ю��s�dC 2çWU/bAGZ�B{�2E�Ī9�7~J�g�_�l�E +���Q;��M6���N�8��1�k�����=�nE{5����v�a{��k�ӠT{(�e�s5>d����g��d�h�z�^`_���o����Ͻw�5|�̳���{Sc���	�s�������b9���L5n�3zƍ�<�0ʖWB���`ֱ1�b#��"��z�R�b1TԊ��C�3O4������Q�s�kT��a�dE@�3�i��T��ؾ��һ��lmYE��� 4��|�+�H�#`�nG�w>tn��M햊��?g�AS�X���:ܫQK�̓V�W5���]���
�A�;�|R�n��1���.�Cr޲�)
`��D��� nC�$Qs�C5C��8��E�~��رI�V�p��6���
o�h٤ߥ��f���xH�B_���R\�@+�w��
�0�
�CMP?X�|�˶�.m��Yg������V��G�K�گ�@U�~��C�H������F����߭�c�H�T��ut��8`&O�/�ɸ"����Y��6�Dch&-�.4�U.%�9M�������r��=H�z����3���_�����xjΖ�:$��*5�&����U��T��Vڋu.��}x�i<j���Cz
�]e̩	���#���S�����M\E��׷�'ǲ���s��,��*��G��UҜn�]�u�R;���뎁���������*��Z��Ճ��3��gh����mXw��n�A{��`������-UȘ��^@�X 7=�q��d�w�go�VaL�H�C��S���b�^��I�C5؏������e|)Fҧ��r�}o�C���kud�����enJT~�qO�)	S�B�Ma�9�[���a%�
˙cc���q���6�,�O]���x�w|m:��.�r{`��YcoQ썗(<��Y�zlYD���S��Q-�1�e���)�j2��|/�!�b7p�Y���*�u��.�w�}�DL4v� #��o+���s��tCXWw��IS���Pe+�_vB�\Zp��K�b7��BZ���U_�f�.��`��<�ɱ��xy.������f��K��o��d���Q]z�h�7��
�n����)��a��vȫ7�Y��y��ՙ��L���P4ۤ{Ͷ��5Ǟ�S��X�!�b��X�Х�.[S@��Y�-+�Z�j��i�bΖ>B�#���9T*�����֐�?+�,x�����\5���~c������0��Hr"��
J��Jh�`\�$����\�>Hq��>����wO�"�P0w�^��ۍxY��)�3�&h�{��oZ"N�H �Fk?}>��r�HN:m#]b&j��1�x�	v]��p�VS��F�M�����8X��FeHƷ��`�O;����^��7���9�SǺK�9�<�xy���nηc�2;�� �l_�tQ�썭Ak�؛Z!-������TԆ�� �6ȉ�O�.��	�\�{������M��s�5mn�)MI�8T�g����?'��!���u-��X�����v��*�U���Rd#�EZ	�ӣ��E\V85�f�lj�j"�yBK6Huaz����
�C\��5����6G��l��s�r����/ 7�'��H���Ɣ��#{��kK��^0j6��*nU<5�� 9?n[xF�G�k%���(��(��$* rg���/�Y���<�}2�R+5��f���\��ȗO^�\zkn���}M#'��T�r� �
Q������T��*�Dщ ��mB,�R޼�M���z�����hJ�()�,�FR4��gy�CK���M���kR�/�������?��}_�&��4�2��6��������[-���j��>����oQ*���F�3�])�,�|`�LF�� Oc�f�zX��-�3"�'���P��@�针�/6����D��8)�1�!a���a��an)��%|����t��
1$dT���^H,!�PI0ur=�[�і��8��%�� |�W2ii�z�� $%mn=r:��qP�4(�ܚ"}��tE�_����T0�=Ʊ������<u$,ǋ���� .��z��׫�r�ϣzB�(�USc��<ȶT�F�O���9׆5)�B�[lam%�:u��<�@�{A�d@��kJ]�c��Ñi�U�=Z*���n)����!�%��8E7et.-YPn�a�U�G>��4}��h�+�]9�l�{�S$=z�����ۣ��Q^g���% K���r���\��-8����g/��]��x���NTn%�D̯r�L���{��Ҕ�[����'�:%D^N���b#�~�2�����C%l q���T��-d�$L�8�����*Dӥ��(�g���\��&�J"W��K�B����9&���
��?�~�Cm�'i������]�e&�]ʣ�m���j��
�XUeI�o��"g� �I���S�S9k��1uٚ鈾�,��i8N�U���҆���<�BC�Y�Y�xҳ��E��M���i���B�~&�J�%�1��݊v�^��Y������-�J�ՓT�c�Q�4O�ʮ[��_��ֺ/f�ɦ����P��'[��&�8�������0�"Gp���ۏ��P,�������y��T������]�FO;��q�͋��T�^~�����ѹ>��H�Lo�vO�\�"������bRs�\AZ�/jF[�C1��vG~zT�O�{��������)����Skm��A�Uh��m�6�duA���\�jJ�Ĕ�h�m���[ؾ�є�hQ�99�E�<����[N��H�#�TP���fY��Z�O�l)+��8Do��gQ;�������d�k���  _�Po"�xxX������E�������>?1����z�>�IpB������w@/���� ���"*[����ŭ�~{E��O�h�C�p�C��[[q��J�6�J�