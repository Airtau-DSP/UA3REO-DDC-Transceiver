
module debug2 (
	probe);	

	input	[13:0]	probe;
endmodule
