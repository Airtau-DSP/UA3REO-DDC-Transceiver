
module DEBUG_Q_TX (
	probe);	

	input	[15:0]	probe;
endmodule
