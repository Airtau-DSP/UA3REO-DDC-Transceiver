��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k*(\&��Y���z��;����1~;ó�!E7+ Uߟ �v��M�a�v���]�P9�Hq��;��p3u*���)a����9�w��mY(���Fu���u8G\��:��^��_eb��.ڄ�f��h��(J���?�G����-��vP���y��+c�Y�����=q��%�h*���h�Z^��=3���f����8��@@ޕ��`́�޻��=7*�K��vn�餤6��
�}����4�p'Ĺ�3h�x�N�P朓�[Cor�%/a靉7]|��d�%��������4�,�8mz=��X+>'����\�Y�����F��������.�O|�'���n?&��͘T���hGS��'��\�����0`����S�dn�.iM���Ц�6���"��^ӓZ� ������a��SxP�v�q�U+:ӄ�Cnc���1~�ETHS�L�I���Fm�Tnj�F�(Qқw�0z����[y�c
O�U/���,�g��^H�0�?&���zj��G�����ɔ�bAl�9~G��ڈ��'�)2T���9�h)�M
�|}����&�,ǜ_8���NS�y��sG���.�n炕�����*�9���c(��ً�"!�������FmK��D���pQ�=�th�v�]Ll',E������9AcL[���2����֌�-�̵ā�녶�·���y�˦E����.�R�F �aq�>��Id6W4�X��)������&%3�Z�c]"z�t�W橻�R�~����LNȞ�D�hݘJ�����
�)�{R�H^(l:rkp�C����X����2O�e��x�M�� ��M�H�1�*��ֹu�4#�e��&0E���� ��XOz{3��������Y��t1Q�O�lG?-�r��@�w:������
�����\�J��S'���n`4�*E ��<6�+��<T
E�`����V�GPR�ԟ|�
�)šy��'�ԞZ�Q8#�G�HC���P��3î8�-���x�z��9R}�ep���X�*}*�D�߻�������?U�SWSkV��u�ZV��p"�9�T���L#�$�t5,EBD��􊉽<�"M�t���1D�^��������v��Ҏ)�Zf�e��*>S��Y���	~����u���A�\�~��t��x	�������JJV���S�k�B�����pm��|�E5��.�N݀)!��� ���;�G��-A����1�7��#�W�#�?�����9�DU����&��[�GtQ3?}X�{�	J�m/2��TiU�O<���leh��Z�6���Ֆ�{n��0V����,\��aM�,p���]��/+%�_3��wi
��h��I1��[�h8&g7m���l��-������ŚcG�8Gf���I����͚bŤ9P����o�M��,��9
g_�� <Jnq�B���&c"�<zr!��JŮ�Y �Ze�\&�M�P��(�w�j���0ӂ��j����L��nc���Nb>��~��O>�5�n�����sZD�+J>�v��!��!O�����Z7���n������Uw�f"l������wyHH����<jb�2�F	)��H��ub�k��e7i�zń喘��`�� P�$FC3����3��d(VGJPfե�U��?��	:�aX^Ѓ�\�s�v_�7�:ʞ����B�x��t��|�@�3�`�u����:S�.�6��}@�t��s�-[���3�pe�U�T3U�$�lQ4�w���`�c��8~�����~��o�5 t�@�u��/��2m�]qc�
�ժ�|�'�Vޙzv�1��*�K&;ȟ�m�.\S��`��)�H9����e��i)�T���V3�!�N�š�|o�>���=`ȳ��F�Q�8Od�n^ef����,�a;x����P��[�Ȫ��,ͮ����o�liR\�2�~�����\�u�BB%!/�?q�߷���?� ��4W}���E�+������&���O��"3���4B��|G*UUo�|^� @="m��%�ppeĚ�N�@9kRc[�~]$�2���{�ida��w"��u
*c�RB�2�!=���B������jL U�>�����)6�V�f�w]/�C+�B�n!�vg�EJ[+�q=����)\�a�qH�sgO,UC�$��j(�C��Ǆ�71���%^t�4\d��M��y�H~�8m� LZȮxʆ��tIƀ�y(����M�s,O���[����4�{��s��;�ޟ~aN��HZ�4n ���{O�T-g1ڗ��y�yΞ�eq��Ŋ��������\���p�Dm�p�Hg!L�]�y)}@�p���}�l8�	�R{�4S��M^��*.WW�n�.�
Μ��)�a���|�S��1{�0cz�b�c�RۄR-Y�v&ۙ-���ƚ]R�Pž>���'�x�����9�_CB^]�@�3�`!O΂!�h�>�w�y��\/���5ޏ+�R�x�#=�d���=gත|gW����E'���^Uh���g��:��gX�B�:I�&��3���˜s�-{�w
[���%2�Mt�g7��������9K�Įλl�m�
g�-T~��qV�X�}~f�Ε���k�_%Zʎgg�bY����	؎+rD������.��H �Ǭ�9dCq5~W�fJ\A`� ��sɺ^���ѫ��\à��y<b˩ "�^��ToHb�a�N����"(�A$iQ�ɫM{���b.f8Ӛ�.9ˉ^�aW@q��H^��4���PU���ŷ�c�]漤�Z[X��Djv�Y��<������1��k��?�L=I^рR`!ؽ6tz?W��?#��L�rgsX�wd�KL�Z�/ڶ
\�'^������F���*��z��	Q��)���^Ls�4�Y�:gC��ԑ����Wö�>#�c)�@�ϬG��V�s�8��j������8ef9M����>����Շ:��mEBh8�}=-x���e���8N�`�t���ñ�)�����I�S� �����A�'�C~,R.�:.���ɮp������G$���o�{��%�;pA�}�Ɲx}{�� �!cl'V�p���3Ӝ;W�V͕���H7��5Bn0K@��b����gc»�3���o^����$�s�"�H ����`y6���`�or#s#�����YJ�f��У�\if:3pAD�.��zS5?~���9�f2�^EE��Ö��mI�y�Hz��st��9EA��C4�I�ʣ�?+����B�F+��|�E���3��1k�5�,���jJ��̦6�6��m���R���ޕ��h{��ʐW��ۻ���a����r-����E҂eQ8�R߾�l�g�=AH� .��p����Nn�5���|ɠ�Zgsu{���~��Jm�
�a)�ɇs�@�V��j�7i%���}|Jko����R���V.�9����`j��6�[��E��Es0�3�ˬ'<r�Rߔ��E���xz���ʞJ�X��+N�\G�Z�{dU���ʝt��E�M(s����h�ys4� �﫸�A˾���I�KY;���f����3P����z��ѿ�� b�ٙ�<Q6��0���3���%�+6Ž�:穂��[�	�A���.�i�-�Z���r��~\�W��%T"Q�9��D�C1��}fb��z��A>���4����%%Iٚ���瓩z��>{="DB�.�bP�rU�5z�H\�#
�!�-�(�'U�2�i��|��B�� �B�c��둪\J�X�W�O���\1�I���c�Z��i�}��;�,<�[a��<풽�̇'?Y^�
#�����b���z��� g-����d�D�,�Q�Y�]֖x=�d�.߈���#�R�y������]Ѷb����3>4� %�3�F��q�Vދ���qa�~�u��r�q�uV�=1yON��[�_��T��&��T]����ϝ%�|�R�BJ�ւ��l[��S��Nf4���2i�i�-�/��0 4O >u ���-!붡�n2	�d5����	��,�#`�����G_�$���:V9��?OK�=����x�I���BKJ�,�7��,7빒�f�=�i+m%��Z�7��D�*��w�M�1lh.(5�'%n�����.�k���ҟ��0�s̏^mrbw���ԑK�����("�8�24ٕCVH�\H��;��AgR����e&�#�"�ʫ���tV���ęs���
J7��{e��TuA��6�/�1(��.��(�^~��Y��f4�=����z{����g{��@z���	�V��@�u��ܽ2�q�tɗ�>W�#'��o���=�9#JD�&a����n=|���E���>"��1�gݦUz���3���_3Xj��!hf��ݣ@M�'ި�:�n�O�¶
����]Қ�}V@��� �d́��O�y��,b�<����F�v�f��|�E��<|ﭛ���}��?��B'��@+5�)�G0�Q�t\�(�6�%��	ifP���=#*��.�~Y��P�]l<�I�0�Z9NV��./;y�MWU�|����N8��_����9j8� ^�g}�����V�ɲ�wEa1\��rj�9:4x�����Q�K}�//�;���IԹejg	u�0ͷ�/x��_O�XvE��dE�\X�v��}����� �:�Ƒ�[&�̞S�wR��Bt�@ʚ��HT�@�{�+�};\�I+��iX&`��g��n�>��
����6iq���8�P��N���ħ�\�}MHX�;>��lL��t�f֟�u��I��|���ִčp:�%�2�-{��Z(�ğ,~��Z��T')Qz� ��!�!A�*8�a���p���2�w���t���hSs���QK\Y��V��fs9������!���mU�Z�M{^��h�Yb� ��¶�s
Հ�-�%�k�m`�bX��f���π�z��/�-����.�ĝ�y��|��V�{�i�.Q��ͥlӯ^X9R��l�	z��8��u�(�$>��G*�0N�b�B��OR3z=�i�匋�;�������g쐉g��깧��~"��[?\˼|>���nyoo��T�^�gu�ϐ`
��x��D�Φ���^o*����̛�0l��^�l��?gD@� ������LMӴN�2D�p�t��|��_H^B�R�w��>���2G�h���vŽ��)`e�S���qpP��-�]����%�%�W�P�z7Ȉ���X�~��o�L���m��3
�&NJ�A0(U�/65ҁ�f揃�������5R��%�w�*���n�_��M/�HSН6�-fi�v�7O� M��^�.�����ӒE��.�g�$�m���
�m���N��[/�u�%p9�*N��$��/E[�������)Ǧ�M�2$l���4�����,��,Ӽkw����D{��'_�p��~p���������y����*��J�1�CF)I=H�y$���ٺ����,ߙp��ap[S*7�hߥ�Q����;װ�d��0�X��h8ZD緭@�u�s}�{@Xd����J}�?�