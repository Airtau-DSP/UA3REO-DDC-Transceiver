
module DEBUG_I_TX (
	probe);	

	input	[15:0]	probe;
endmodule
