��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�����S�%l2���t�y���O�wb�Rv�m�����'�lٷ���
?L�����*�FI��j��-�j {�G���L��#��x�$�\�ի�yj��2ݸ�=�4{�}W��
-�[[k��!&�m�ߤK�i	�E7ǉB���g�iؖ��X)�UhX�]����FP���6�ctU������I��$OF�����=�i����Ya�e./���9O<�����e}��FA�9���:'�)��͂�k���8�[G����zTP�t0᪱\�/ɑ�3렭Y�P���	�&�<ɚ��2��T/����_�?��{1`)}*��e�2��Hwsh�"��U�Y�,�s��&�����m��E?�+�
��rLY��JQ�)љR������}a4բ�e��
�U�D�E^�|�~���`��M�Q-��mb� �T�f�Eu�S�:x�e9�����xS~���հ���%�����(���;��y@pXδ�j
����Rx_tPH�vD�\Z@w������?K�(hm�
��#Ҩ���,~��xz����Y�UAQx�,��̮�����G#.8=ښ �X(�����C��%�\��R>b�������R�6}*���N���8|9����=U!�D�c�D��I/�,�<|)Zy
�~(�({|R%9�F�8��fT�o�).Z$�(�����gB��v_���/������GF�~�Xױ��K/��AZC{�K,1xM~�8��F��ź%QQ�ɬQMvZ�L	�K¬~����)/�GO��G`'���U*�Ƨ�y $1���<'��.�k�eV�06 s!�6Ͱa[�V�ٺ��_s��t�f�`o��x����D� �n^�H/̸x=��Oh\ւ؇y���캉��P�)y-.8p$KwѾ7�V�3v%���KP��s����OV��T�lP��@����ʯ�G������s�"|�"�꯾cJ��x��u��e��E.�
���~��I RCJ�g����t��D�#g����E$��Hz�i��15��($u3<D{^�z{�MgY�z�o����rz�;�#���͞��|��,�'O����-�y>�E
k�eIQs�������mU-�P����gYM�"����u�P(��1>��-� ?a��l�@5�Ѹ5]�c�<���6i��HF�[��Ѱ���"e�M
���aI������##�U�b�bu�6+����5�W��ko��2rλI�z��k}p����d��`�Yb*�F�O_��c�ya	��O�	�5��%��WVL#�s��L
I"D���ø@rx�z�/��AO�� �Ѯؔ�FȬ~�O(��U�+���X�<f��Y+¬�L��ztCW��wQ�k9���N;?�D��R��|��:�yNی+�.�~K�7v�K�f�,��(���7939�@i��F"I��j��NY���d}�'Ӗ�ʢ���
qN)vo�� X5h�K.tcW d�����]?+�o�M������
�y�T���$^o�:��	�[�1܌\	���Jh!�^˥X�G6����^Ԑ��ݷ%%@��t	�6o8س���=���O�v��N�&�� .4����M����
��7Y�CB�W�!��"A��W�}�*�"<+�J:}���D�ϗ��xԱS��c�AyR����+���Oi��c�����W&� 9��X�Oow(l�@�}8IZ(G�������x;�EJ��P.�D���H9���%�ר�(Z(�Mҳ�6���>�W;/P)�.p�hLF���lj���K@Wϧ�N���t�E��k��0Ճ��p�<���s�9]~�F�j��-�Wp��K���"Fe5I�A�0��g��Fv�ǽg����|4[���2�L8�/��D�>e�{O�q7��ƴ����`�g���g0�a�!���W�~���ᱞ�E��)���R��.�@x9�5�ܩ�~�ɽ��InY��u���ɛ,�@�V��$>�U2Du�:��2��M.d��#�.fF�	�*ʲ���߱ohe���ԅԛ<�g�Ǻ_ۧS�ъ�Z�V[؇T��ZP�"q2o�[����R#㗂��Z�.j��I�i_�В�ɧ�sM�f�Rv�\�,�=!=׼�s���A <eD��&��tRێև��xE��p��et�"<����N���F�������?_�l@�m)7���K3��v��\\;xcDr=Qh8�jRD�Q����s5�w�<e�I��*m��XX?"���4���HD�w�,�A|�j)�r	�ڗt��D�X��/�È�Iú�qGk�EU��]8�UoS����ĝ6�2��.���(�
�?R���#��fǽ�:
7�P���V7�};��Qc��7	��#���K9�U�P�~z������+�GR�����:K����[dm�j�V,(����ǉ"����.H�c�	����K�y�3i��˦�ѻ�x�d�u�#!1�N,}<#m�I���
�a�����I��q}R�5�ׯ��_�<�NrLpw�	�6��(ι�s�?�>�la`�a}燑��M kcY.���-�*��U�N8�j/�H��m�L��bE�!i�����}Aʿ��e�sؼlF-�s�uv�İ(s�#��FSG�noխ,�φsx�D@BK��G����!ah�}f�ڼR���d��(}�VaU�$�X�}7ʀ og�� ���RLgF#�ivų��
��{x������]hj� q]�x��;��ъ3���da��Uw�+5�xAM�K5jF_��TA�\���b�6%����(�Cc�QZ�\���i��G�P��9�F-���SM�a"*J=�	Й|6�n�j�#;W8������"���+��CGz+1Г��Գ�����Z!y�� ��H���n��:�G�!$�&��/�1��i�m �@�0^PW�`�:����IC>���?ë�r����߾�в�]��<�r&RC�sB�m,���ǰ�Mj���b��q*��yʯ%i]s]��) @�R�ICή&z�7�s�	�����W��T��ǍDҲPo��Ç�<��o$�}��WE�:q��oѿS��`:b���"bL���P�V��	p�)T<�B�3*R�2�<��U����VyQwF�$C��ћ�u�ۋ�.��g' 6��}��$����UK�u���v�Hs�!X� A@rՕ��o�np�&:m�P}��Y>���2���Z4�P�Oa'Yf��X?�Ə�0�����#��?$�-�R,UC�QJ֍��m佔r�7�ʪĩ3�!����O{{|�w��jY�=D���Gj.3��T`�HS@^g�	}gpf��G�1�hs�6�0��޲�/�[㵔�j�ۍ%T�Tܹ�c�I0Ԏ�$�C�EH�1D��i]���F5ü��9Ā7�(O ��(�^��Fx�Θ�"~+�S�o2�;���ߝ�������<����w)��J��%�j���8��Z���\�pI��Sk�٠��DS���ò���9���Dz�2�����,�T_Tˎ]��Z`�b��%L)���+������VnU.C?�������ܟ�R�Y�<�)��B-���;��1[�~ N�X�B��3��>�bY0�N�8񒈼ӳٕ	ϑ��o��[4�0k�=� v��i)�4��ΖN�̧�[���A�ذ�uL�|S`U~�����"0���*�G��,v����1�T/�cm����o5ꍄI�Y��k��TT��)���Τ���{1I�t��+C��k����łO��O%�M���s^< ��R�C�A<���Yd�V���:�.	"�!"N��5���N�Htf�����"T�֚���e1?sv���T����3C�	V`�����M�)�
,"7�[s*�����,������aȠ�bENW�ї���k�֛ٞg�OQ�Gk�DN*�d҄��m����vt<�!�}���r��Lo�E���/CV�Bu�����M}77!L�.RB	��75�/��gn4�nש��ka����p}*��_i�3:8 )��-���NC�Y\%��@�fK��8I��B�Ҹ8�g���}��؍l�u����I��d�$����T�O+����e��	��_v	�jy�f���i�� w��!��n)�s����\+ahݰY�O�!��
�ܑ��p�Wή8�0[��G�u)X��<�5���$0�b����mQ�j;�<��X�['��:	PSx�#�|2$tB.