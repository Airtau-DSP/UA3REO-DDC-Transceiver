
module DEBUG_Q_RX (
	probe);	

	input	[15:0]	probe;
endmodule
