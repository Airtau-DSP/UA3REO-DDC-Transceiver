��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k*(\&��Y׸4o ��B�w�P q�D���(=_jq����o��N.Ұ��(n�L2���CB��G�1a�-͛�ı�@~-�>*QP�����]1㽖�� {��gw�lS2�$���(ǫ�!�^\P�؁����K�*� �V��EE����y.g�#�f�#�e������6�7�{d�Z�#`��K������L��{���c�
2o�a��׸�g(ݩE`@��K��c�)/��wBL�P�`C|[�2��ӽ�f�A��㐟��i��g�ӄPwj�ےaN�lK�W�N�z�o�YJj�5���x����FQQ��ޯh��ӡ��B��2�Ϩ�-���wV��s�4���B�~��bel��=u'�Ա:�0�08C�ٔPB�G�p�߈\�l��Y����u�����O�Ƃg�P|���6q߄��@��ɊH�q���c�#G�6,�gϚ|Kty��&v��x��_T��l�R�	�\�T�OG*��]�ܘ]b�b�o�
k��
o�l��*q#�'M�F�����!��U�^��Z��$]b��d���FS:u
����_�<p��n/wWg�!���b:��K�#�u��Ė��-X��7m����Ǖ�f�̝�����DU�}S7ZLÏ�ZQ�4x�Ʃ�f��X��L��	���S�s�U�I�y�j������d��N�6�ے`E�q&S�3�:��t>h�[?RŎ�T���S+���8�G�(�%d�ʹ5;SJV*y~�"�*ɋ����b�|�rˆ��/ĩ�����E6�2��{h�
O�����D��� Q�f��wlL��u)�q	]��+J^�Q҅Z���?�*5U-���E�^"2R��믙?����.o�+>�~>��L����#L���?)�~�[�2�zUA9W]K^��#�Xb"���wE��u���<u�Ρ�$�Rz��=ߍ`뿐*��$�ʔ/̪h�z�{ˍ��iU��$�A����Ɔ��q|��h�8*z���NsK���Zi��LD�6oP7\�a�#�<p������<ӎ��@�X�=�WA�u쿢���� 13���Ilv�x���0"=��3��IG�����-��u^�R[H�7����:�_mˇ��
�g��U�:�a�BhA
�x�+���s����
��*��8�h4b�Ճ�u�*?��B�k��XE�'���/u#�O7\�$���vw�]ֽT���_`J,�M�	H5"�~`�@B�e_kt9���w�a��b,U�F��ED�<�0c�w��@��5�NEXm�g207��]���x?���$�=��eZ����]�6S��7���w�f����*���i�"[��.�i_����T�϶H��Ӆ����K��	p������x��8>�vI�����5�C��m���y.��ϧ���L������?t�\�VӨ����4}ԭ�q���ϬYX/�%�*��M��o!
ۑ|+�9�<�r�@�msy�hyR+����b�'ZY���R���0m!�NNVh�O.�dF2� S�Z=��ާ�m�!��Sv��(��6��-A�Ja�T�d�[��������(��~�M7�g��&BԬK��.W�Iʔd�F��3���U��|}��L��Q@D|��V��}ΝLtw��tE\��*��/�^�^�?�O�@܁����6!��C�D�|ﹼ(���5����G0m.}^� ��$
R�5
�,N�m�2���^��x�����M��5����þ��l�2���qÈ�e򎬘����,nn�G�h6v�_?�^��ԑ/z?��F�e�r�N�Ql�o|�bV�Ěa"{�9xD�m��~��B42�����S�J��n��/Aե�g���D�i� 1�|>_�����~�Kc3�66�K�����dP4=T.�Ƿ �&͂PKV��WR�е��kg�a��܍��ur���/s���m����=%���V�����M��]$��>-�'��R���k�o�y���&�~��o?��o,�J�G`�;l8�C����tw�l��獊����pG�����r�B����k���(��x�Rw1����F��|�n��;+7�#�ݟ�G�#�h릎�1+�i�^Z���l�IX��.�κ�_q~A��?��HަKO���ooT�E*l�[=z�Cτ!`���s����,�Ϲ�������$Y<I Y/@�NH�2�	(�	�z��t���S��VZ�L	�JWQ���(w�sa1
��ŵ(غ<�p��I"Dب�E \�}2�o��*,�v^�?��
h7	�)6e�w4TN�$$2��}h����(�(��KXx��!���ǘ��;��F�AW���W���
�a�5?��ɦ<�
�:l�u���fO���J�lC�D�h-�������N���E8gq�C�u	g;m'ЄsZ`�K�qPb~�-���$��"H���z�Pn��C���{>�� rA̍cV_T^Y��y� ���]M�7>��"�x�;���qr�K*����`��i�1�0d��cpX.c
nd�j/;VF6�3�<3ؖ��\�uv��s�Ҁ�l���9����?��f,��Ψ�.[�$"�N:I���8�����#���w��#	+���}�>�~`�tww���WS)���P��yC�������)�>�Q�l/6����*ȥ��5Oݝ�^k�o)�Ry8� �=���N��1������F�c�&&U�;�p�m�F��?$�w9�U�ݕ����Bpy����܏�����aV�d�^��\ �ϒ�8@�CJ���d��B��������BR�Jf��%��6��y��g�c�E)�