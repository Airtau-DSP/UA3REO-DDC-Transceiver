��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���'�ʞ�~|�A`�U���k�,�ܻ�zc����9z�n#�?Ff��w�Ϯ��^�����[�0�=3i̬�S��
5N���-)�[IN. �b5
��N��@<�"܄Q��X�q�E��?���^�Fǈ��������0�X�(�`�*�y���B�Ą�-A�Ua�D�I��q#�E�x�!oӔc�o��SA3��b���\����a{��S�e\����.�K����\��J5l|��r�2�/�.S�aΎ���T�����������~E�4e��7V�y�^�F��{�yV��G��1;��,`[դޙU���G���ੵ�����
�ЦT�l����m�g�uH�8��'�}������U�*�X�-�ǋXԲ�������O�' ¢�uPQ!Me �Pp�,�02�aW���S����0���S�#��D�Z�#�s%@6�O�u	�q>\
i��[��'�3�� 1�����7���,�u��P�8��i�;��~�\�����6j�yɢqù~S��=���Nz������V9�8#�9�#)����oycnD=�]~�W����ȗ�x�"�s����*)l�j,@�.�Z�*̐X���gX���n�H �@%������߲%Q�1	��;KZ�x��0c���Պ=�Ӻ�Av�.��?��qU%���1����Wf�P������0����:|$+<}���ݕE�Ks3L�)3�B�y��o���u��{�-8�S�F$xf엽/}l���{R.bs��ҝv�?)0�W�0�f'�0�m	��6����.��z�S#����@M=��t�XH����b���:�.��\u?¡�s(`��.�ɢx�/�:[Խn��Bzq����,�>ҽ��1��<�A�@��7�挍��tW{%���,He^^�]�o�p���G��6�S��X}@bBE7ǝ�<_�K�)�e��ℓ�0��=��#d�$_�T�� 1��t��N��l|������X���l�)�7�-+��ΜK2Б�v�u�kK'xA7L4��ӵ��Q�`lJ�O����GZ}Or#�BF�1��SFr+��kJ��B�.$!+��t7������XsŃ܀4�6;o���;
�ʊ�S��et«W�6���ϒ] �B��A!D�h���I�f���P�xn�H?��~��3�ȳ��\xȳ�(�3�NyrY�<mL�c��4��nC�e��+z��gJ��FJ�/��{��deI�+Iy����)6gvp�;\{> �dOꍟt0�nV[$$Ĵֈp����?�Ir�2�,:~�;��-�;��fg�/VK�>Zv�'�r-v��i�u7����#՚��﹖�I��퀯)��C����[x�ٞ[O
�=��h���&���6�+�*�w$��)Y�R��y��i �CV��2E���ʃ����<���#�.�:�~E���>B�.�L��A����\1�N����x�h��)�Q->��;Ý����ސ1����� �S�}���A�^a�wW�/+H�=�U6K߬�hm�*�_�{�A�w:7}�l+j��F"M�럂���D�M���J|錠��(��YIh͙j��AՅ�!����~�4����ׄ�%���Z�q�����ё�[W>1��Dw߆�S�Jo^ʮU����M�09�mi�c$' �0�(鉀;�ǆ�փ1X�*&D4iJ�Ѝ�w&�{�9b,�oe*��j�^�a?j=_��2O"�&��*ސ��[\�&6�%��{��]Pj��8�LZ�����S,1�4��iJ����PR�,1�����ukѓ_�-a��P�y!�NvުB"ˢj�P��x����Ցʌ@..2�)0g���j���z�� K��wD=�?$i��Se���k�P�(����4���$��`�=�uA
�A��V�I�;����P)��F���5���)�G��m�m��.S�̍h��F!Ҟ�GӤl�ݿ��̎������Xo"*'���s�{Ղ$m-�� �nߞ]��۔�Y�Μ�c5}�jg�5����r���#G%p�������k
O-�ִF|�I�3�}K��䒥�C5j��m���m`��\'�Ю:	����V��h9�(	f� #O�z�/�I��#L��لv��.��Rg�6�
�]�G�kJū�
b03*4�i��`��5��s/Fﲁ�q�����eZ����n�����~��U�lE�"��8��W��T�n�-�3]�\�c����2�=�"������C'�l׽���ؔc�40�q��LB�� ��6L�o�,O�\�m��5��`xRt�d��f�a*��r��+���W7����?���c	����Q��+�vƲ�z���~����h���0.�j��+vt�˨ނ�}0�i����`��jG#���+W����Ϲْ_eZq��W%��	��q��{��ጰ+�P�ك�Q��
w��DU��Q�����d����	sU�(���mc��z�a��?��8������F|wgU�C�)/xɣE�r��;w\��ar���؞���[-���^���o�f�̼�5$Zl@�!9���`��^�-�s�@���fqh���A&sq�R����u�)x�$d�R��~��\�KZ҉ۍ���dBUm�Vy���.�Tri�������iV�����\5�h�=��r-��p+[B�w!�,���"�}4�^-4J��v����7�cp�o� 6I��ǑtſݩN�~Z*0���7Cb<
nf��t�^�R����6�~��"lk���\����]�h�`�0�i�%�A0+���ٕ"l��B#���e��i��8�0w~������w[CJ�8i�����өq�jF���л��}�F"�(=98���%W� .Q}��&er_<�aڣϽ��!�����y/�gE��*+�J̷ݞ��Dc���Hz�4u!tD�JKm��� �����RG��jȑ����,�L�tZ4/u��&�C�D�W\�[�v+���-)�ݧ��QgG4�n��n�&.^~�jD��~!�pr�k��J��ِ�A	���(j�Kӥ�UEp�v��n,��'����~v�V!�\y��(�`��dj�~���\F�hW��^Qz\@��M2{�h<^�%#I��J;��}����h y[��>�WM»�����S�z_L2�ZQLd�u�]FK�p�K���C�R9��WD���gi��Hm���p���S�s�|��[���� �Ds���-]���H�B5@��6�LR{�Ew.W��s�ry��X�O���s�	��S��'볂�gk&[U[=�b�:�fk�S�D@�|
��/�;)U`XC>�{_ �`��c������,����+�@@Me���&v�y�}�"���+���_7�\"��Xlܢ%���h�v���q˂�W`�x2C+K�'q���RL��1k�zX_���sz>�\�-�s�����^Ⴣ�@R��v`�{�b�х%R����4�Xܣ��Qp$b�1����I
&��fX�.�[���Q�'�+���^��Y�>� �Y�Ġo�wwQj��Y�#f{x�L�è�M6,"v�����`u���}2�>K����&NO��
�!�J;:<8#�ߺ�I�|����/�՞�ʑx?� QF�|?����!�;���F�6|`�%�'�9)������͹����:A�� �=�G�3��b���a�F,��o�;p����FnsP0k6I�T
��#P|6�N��ٙ{���p �������_	�u6v�@��xk��ä�0&�_$���/��������E���Ln"��K�&m_��x
�RO:�q�B͏ȯ�2{�!t�9ڸ��_��2U���]�L���X8����� �����!�z����m
"��Y�wҲ��Kvyީ6�{4����h'0M��qn��g�Aϰ$,�^!�\��cp���*�"����L�Q��c�1�B���Q����6=*��]���57����HEu�0�A��!��|6�@���`���+ANt��恰���l�E��F���Z\ͼȂ��AuҖ��sؔ/0!`@"G�!���v���	Q׭����d�Wz�ck�B~4Xz?y��uL�oz4A��n٥PH�%)��-��F���Y��SO���͕W����fc�6��L���׼�Xg+ˢh<����?�`���~�d8���0�7��b��XzQ��e��8�ׄ�����ٗ���I�I-~���Y��p��C�]�,/m�:$�T2T��q�E�}j���{�����k�}�_�R����eP(9�$������މ,�P��5/u�r�λ����%Jr$�^A�j��eEIW0vɶ�br��8���j�n�w�ƳYB�)B�(6�He���ϳ�	�HJK�h:B�J_��6�y�8����;��9%'�����'���7>���Beމ2s�o�j$�d ����
�:BB�rKw�\��k{֐���cNk�N�J.Ifk��+��;���+`?��MѮ�k�%g�~�d�WP�O��D���4g��S4�3]��	��#y8��MЬk��Şn���i��o�A0�Ui�|�r�4��w��^e?ϧf�Z�,�x��G���<��O��剥5�Sv~���L�K�4%���b��1O�#nJU��ՠ�U)���Tj��d��n�`<�b9���a5EX'�c���E�����4�G;�I/�#��+�s������X��
�i�i��L>�.)^�q�J�����A����ą��P�F`�v���i��X��,6�:ܘ���u+J�%��O� qɢ'}b!@B�\����(��q�I�F8�&���o	�ghߵ�$Q�* P����pjO����v���M`K�6�1����?ں��(v��W��gf�'3��&`��$,�P9�j~��3�$�h�!��R��2{����\aϧd%w_"���
^3�2�M��}۬Ă��P����PS���qnO����N֤ۨ������)+(�x�-�/P��T�AZ����U�No.�1z��Э���V囀�4��^���m}���� ��rd�T�ϊ:�ne�|��>d����oR���?N��P���o
�䤭�n:|�yC��/���Y�S����C�u;�q�Ĵ�ri��k�w��Ǭ7M��� � �z��P��2N_���e����\�lu��O�'��#�S*�{$��Ŷ�~)&�{���0).G[�w^�8��᧿����$��J��U'/3c`��zU��,�%��q��}@��V$p��C� J���pp������?���I��dJ��HS�7��P;y?'
 �ElՅIӊ*]�9!�t���1<
��a��&KO�dkE�^���K��T��F�uF_8`2_ ��aS�^B=q$�𳻶�}٬V����N�[�Lf�^>0u�T?t]�o)'*h�[�Hю���'C"�+���Y��#������_�r���%�
 5ӫO\p��c�[�����EQ1���͕���� ���
�u�Ci�ú3�6��M���`�~���-|t�WR������ɕ�UV�p'�WJ�\�I�R������׭F��u�n�l��� b:_Δ'�5��2i �p��,\kSX��"���dILI�Q��tk����u��<�b`A'�l%$q�9N�9�P���
����&��k�7W��O��L�B�ɖ����iT7R([�H�MN����u����WR���7(��P�mV]�%I���v�+a+�[#w�D4��� �f�:t�L�O[AEN䭒��q�.d����E��b;ߩ��MZ��xH��z�Y���K'�.�j3��-�֐ɮW'6e*�l�S��8]��D�����ۥ?���ƙ��C��v�)'k��6���K�J �B���;�;R܇f6Pp��~	q�������Kd�b�b �R���`�,d��d��w�.:���(P�Yڋ�E�ٿo+ ?N����I!u�<`��
8'j�V���kcكzB�y L� }�q��0���l��]<,脜�l��oD��B���Vng����%������V^Q͘�*���ڽ��s��� ֨��D�T��t��=��?��c��h'ReR?c%����u��*�3�wNui�l�蜚�#��A/�}}��0�.�K7�q�@'�[�{5����|�k�`�����.KP��ճvK7���*�1��C��nе���~�}��{�	����J���^C0�����3�̬/�ԍR�ltFg�9�t6P;%P����h2� �1P�9�ۻ0U�<tr���'�d{�$��tɛz4������ݫ������X��p���'��8���%1u0]� 7��X��2��ݟک]�r��AE�86�m�[Y4�Fl��e'�.�F��A+r0@�����Ƙ曼��ͦN"S��;���4=F��i}�j~oD�e�@����M��d����ESЍ� �ۏ��R&�6S��k��