��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����ըf�%�����KRs�x�̊f��r�L��W8͏r��ں�9A�窔*j�D�)��;���F��*�9~�Һ0_h����%)��
3q�9���#?�h���WP��4�pj�)�F��e��R�g���8�y�Qga���܍M��D�/�6&�,��'��.Q��S'8T��Z=�*k��?]���z�)�c/�o0F���r[^���\1.,ɱ']	`M�xd*��V�
 �4�n���3g0�=�́j�3�S���A;ґ�L�yM�Y���&IDߜҡ�3VQ9�W�Th`���hk���~�Q�Y��R�ݦ��`�"+k�	#���:Ƶ ��>|�f�~���9�z�w��BW��_7��S?��jRKK�C��4cǷ��M��&�1����|�nb&�߅
���tq1�Ir���Q/�_#W�V�k�MD�R�����9|�ۧ�S���_�_�ڤ�Ϛ��!°n
#�e����ڨ�|�]a�{�.�֓E�G�j�][��^Hgҷ�j�$�ʞ5ё'±^c��d���T@a�$d��wy �<jZ #�H3�s۸�*�L+9eea�U~���a���F����g�1��R��������h��������3=~ ���կ�U�ա����0Ȥ�cd��$]9j��$����d�K�ڧ	�$N����V߿[�x�̎�In�Q(�Lf}Y�y(af�_�h�̒�����c�I�]�JGR&+=��~o��X�ݪ��uRE��ssZ���o�Vr7�ܲ�q���pz��ܾ���J���W��1�3���>��v���븹 tj�[�s.���'r�ޑ�O\���M� +06fuL��kXW�c���c��n�4� ������%\$�c`����GY5}��K
/s�y~�
�Zg�|�6��U�AuO ��}M �|�;cT�}k��p�s��5�41�y�Q����	|
�F��5����[%�H�P��u���3��
�\����'�s:���D�͛�c�'��?�+�?H�bP�B��v!ٌD��Q5O���Ʊ|�q	 �pg�#ի�ej+r'R� �.��2��x���e��� E���̿�)�$�9�2�!��7�϶]N�i�~��$��~9��2*��y?�}�sX���H�,8�0 �Ke��]�`G�x-�)����S����a�Bk]~5~򂓯�D��>]@�7&������w�;��u��U�ZE�*`c+��y2G�3��Kv��{��{V��~"��rej���P�q/��;u���5����Ve/�*�?f]J˽>mg���km5Y��Ѻ��d��K�$>AP��^J���N���-�B+]�8b�z,���4<���v��<h���@��H'��-��=���A� ����EΔ�{X1:�=xQk�7� �E=�U`��Χ������J�#T@�J�̠�;�k������*i����V#�e��;�8wP�R� �@(�>�2����*�w��x8�>���syd��d����"�I�/���X�v�˂ ��[W��_�-���qRK��r3�W�_�<0	Xv�M^�J0��_0c�d��0�G�y��D@f��ZA��eT-�x O��f�x��:�+V�8n5؞���N��ҿ 푐	�L�����c��s�a,�J;Ǣ���>��Вu��RXJ�����H8�f�@�9)^z �2"��l��
�2:����S�Y��@׷ýH;\��o��Qq?�,�k�.V�P4�IW�V} �vU`��D3�mV������r%V,�v88��W͝�y`��'�#b���Yγ��4Kܞ��/��y��5��*S�T�7eR��a���\��+B��3;�E�����P���w�d[��b�G��?m���>V4�2&r]L�ƱL/�eۧD�T.�0VǍ�j�8oj;k�d���,�$S4#Q]���ty���Pg<���c1����QƒB��Zw(�f����s�j��m76��6�j���ۧ��=���2iҚ�zW@U!��Vm }AVCX�J/��Eqwg�)�0�<�`;�JV�>��j�����:T��Q/(���1��Kr
Ȼ	��z�J�qK�m�b���串�[�Ǹ��9��\Õ�'��^�(uM���-5߳h�}%��V&����:c�l�k%kX'b9I��v�:�i��c-�xb�J{гLE5��9���[�ľ�kb,d������Dw���� ���8I��ɶ��^��Ǌ#~.B�{�ק0!�u��X��J���M�U�s�	�71�������!���V~ɛh��I4�����}-R� _�9f�uS-PQB��X��`��~���=b9RN���5Sf����-�ۨ�4['��C0�5�
}��AEY궧�c���O#���>^<��&�z_���%^b](/������PK,*�v�1��X��g�l�u��x��=	�1�R螟�n�W����Mk�u��QF��m�y�:�'�o�}�*����m�9�Y�Z��k�f7�ս�㲩]�_m����"Ϲ�����T��ԭ#�N����[���<� x
I�3`}3F�Vt�;G�<�s��	��T4�f��9t��L��2� ��"?�K��d��La��Ka]��2���I����e���!�?y�~���dn�>M�Y���s�l��)ʐӫ���Cz)M^��;��-�	����Rx�2 ғ��;4k�ڦ`3�ߞ(��Z��+�f��GX�{dJa�h�:�h-@(bZߥ��1vŔ[���8�(���{?��J��kL4���V�p֨��C8�Y�q�N!�|�1=J�b=�ia���o��< �#l��C?��
3��piB �ݦ
z'�u(�[2b�r��I�9����a�`ֵK/��*�����~��Y��7;�G�|� �P�v�>�%� f/�:�E����0�e� 0�AH������/��^F�%'/���������r�z�����g��	�ϓ3~�z����5L�,8������<SEϲG��aZ�1E��ϭ�F�����կ���<�/噥�k2s�lݫ'�˾nL�5)���N_����zXGH.Ǥ�ƞ��l��	�E�_Y���[��[0�)�r΄ïߎ��2�?X�չ�87�~��5uu�f8�-`�evH�\f��ЏoT��uJ�Z7J�� w5K��2�����"�d�Hr�f�F|7��F�V�f����K?����ʖ������Č_;�%-`�7���l�R�#w`b��>,/�l��u@H]�v����5u�uL^�<��dKZB���a8����xi����Z�\h3�n�M�N���ay��囵1�q�u���O?��%�Z��V���P,yPm��o�F�!�4ˋ1����%��x���}q�:�����{#3������>��1�Y�����1�F+ȘtX��&� \�b�M����G�>hO�D�
�%�G�S�Lw�~v���ܴZ�Q悲"�1v:	�:(�|%(�ą�^�g{(9J�ή��C�]j�Z�/;��	��~��c0�Jk5K��#LVT�⬗L��>9��9��z`(�h?� ��w�C.�dn���yu�z�'���ub��D���P�K�Xܦ�H�;8b�=�iv�f$][ϝ�^�1����f|��[3X:1��|�u�<���ȑ;���d!�l�j*D�'׾�6K�bI&�m^ٚ��P�68pA ��
@�v��K7���k����!��`*�2��c9�DeT����&���ֹ��Mg

�9�N��FЂczr�y��W��}(2dudW0N:�{��=��9�CJ��oV�[�����f���L�=T\�Bɭ�\vl#9��-R(&��+���G����j�.=����W���a$�M�*>�?>��z�'�FlN�6�qO鷵>�@��Z�z�S�/C�ՑB���j��'G�n6 �Y� �X:��m�p�s��o[ȕ�.k��Z�b�U�Ȁ@_ɀ?����ɬ�.�N�"ln���wL��F2���]�b�`�,P����!�Q{*�5�������(	�@�U�����r�����&�-��^��Z0��W�O�z��C�鰷w�C�]�	3�P	�l�D%��;���������b�`��"������:��@-�b���6[�֙�����kVt;7N�G����˸݈h��s�<3�*���d�"�f7��"��][�7cy]����>�L�lZ+��Yd�
��C1-�&?�td�2B��L�)ȏ(�5`PA�-��^��ajv����Oe���E�=l嬵�ߋ
�wxP��-�SN�{�'�e�Dw�(h�8�r/�h�H`�c#5�Ih]��]Ԋ�e��wȹ,�BHR8\Ӡ)�Y�
�r�pĪ���~ß:���r^˝&����8��މ��׆�b�3Ӄ��-�Ѷ��[؎.V�֠זK+3����W�b�6�;��˔V���|�ԃ���Th�:��H`~X�$t�x�W_,�p��)CX����[��'E¦iP��2J��� �1�n���ר2&yA�b�QQ���׭���<�F�ӧ�@��s���Eɢk$���ר��O2�c��q/U8x�J�c��D���鞣�� ����6��f���� �1`"��$�]��>�FO������z�+��;wߚU�V���į�\4s�����6*���']���6k�(h>3�xE�:⮕�T1����Md��DJ
�`t��*4�����8����V7m���$F �$G�70�fH�e(���tb���ֈ��-���d�@)Q�@��:����R��.�R��оfW~AKD��o�	��]M;k_�,�l��dv ��7�����I�76�3N�:j&�b) c@����tq�8�.�5�I���~�QČ�Cv�e���!��&)�+��<g�kW',��hE���.����I�@om�&F��Of��u�����)���8��X���nn�}'�H�
7���s���7�����"z2`>���b�F�\�\H��Ӏ�R�����b�Vm�{�Y��8f6�Ƅw��!=�xwA�`6ZJ�����╢��'�S�I���fY��*i�ڦ�{�x1S[�[9dg�PWyfFȭ�q��*�ɋ���Ht�S���N�B��w�vv �����N?��6�FX�h*�w'C"��mE%�a�����Mෘ���A������ˉa�$����X�^��
liP���e�z �Ph?p�5�z�cI�T}�v.|/��´��qs��h'#}8�	>���Z�Y��ʥ�\Q��3������=�r���}a'����s�i%��\��uF��}���g�	-5b�;C� �(R";H�4�3FG����W�Z�#5���H9A�^6F�p�0���
f3��X�����&�zC����S��N��
���i�SJ��_�q9^��&��!>�N����xQ�N�锻�3Rl^rDM��#_��A'�m�Ӷ+�U��>B[M���}�+����R�|܋��g��,�hw�]?�BAm*�������=�{�s���HgL�-G_��mGٿ+��s=���gB��c�һ��s�:zջI]d���r7T�q6��rQ��f2nZ��#=�F�����Z� ��:
���c>��o&�<�Қ�n��~b�r����-�0��l��hՄS�4��`!wwGjH$I�d�ԡu�S���@��3��%u��7��tTn��l[O��vr�h�j�P������w���;z>(����I���l����1+��i�Z�A�3[?���Ւ~��eu!w�!��u�i��袲]E��{�����3���'��<�x��ƶ�	�{ $�dtIG��ޝ�2WD�����R���y��0���Ε��nnER]�3QΚ�p��[�^�7�<�.���s�=�'8=��-z���-����h<?t��?2J9zV������n��`S��������;��qoU��^�<KJ��3��O��2��K�r�yP��lyfMI\��|0���G+��Z�$*'s=�o�d��'����
��4���!�x�N,W�>������?�o=t�Ыk�S��T���pf�l�v��ˣ��\�^Ә���>��! ��Su��D���O9�IH��S���>��z�L�a�O�܍g(=�޻4V��V
"�A��̶���ƒ���H�9���+�����"aRD9l� �$��l����gg�P4ELD�X�Tk������4.�����j�4BؔH��t��&�_�ګ��Ed�Fa��6�j����]�a&:t&"Cʛ�ɞ���ɴZ�tYlޝ�̲Դ�I�~��w[3wF�+����ӌ'�"EF�e+R��K��ͪѼ	/��	 �Ýu�,@�[��dk'S�M�CJ��d�(�<a��`���=���{�i��É1� �����5��_����@��)쯈[w����k	��`����S�(ۃ1?��t᜼���M��b5a��8�Ⱥ�y�r܊*Yў<��\����7W���i���oۙ��`���ꑁ	��M.��5 �{�k��Z/�SV��&�!���P];��=�ߢ]��LI��G�
�ʠ!l'X{�ڤq�S��m��>-u6�B�X���\C�٤
\FM�X��i��
����#��rP�20�)]L�X�� �IC;�~�8�<��P�b^�����]��a0,���r�=Ɓ�D���K�[@�d�)��=��<����h&��h�d�H��4�4��(hG�W�&��4K?�2X��yMk1�A/��9�����s���ɝWo%��W	�����C=��)fT��`B5�Y#br��uz�����j�
����$y��Pw����c�V���)���L� ����7Z(&��<	�gyx7t�8�l'�ZN�G��׈���7�8d �(�+}6yS��S�y�B�*�*8M�uV�j`�)E��J����mq�phz�T~�ɒ��8U"����2�̵�k����O�)���^Ă�f4�T������EjmM��B]����e��11]��(��x2����A��?��כǲPQE��O	@�0H��X"zk�_p�!��H¹���:����U��!@��A�C�� D\Q"Y
��m*��&�T�[��Gu���\�ߏ��T��	W�nMx�$�݀�T���
m_�!5��8v���>Kx���0���O����k�>���O`�X��8� ���P��>Ft�>��s�B��jt�*dI����k�����T�pN� ?�bɗ@ϖ��e)�kr��/ie:�Z<D;AVI���ֶ���9��t�m�
B9�}7� c�eP�rgO6�6�]b��`��(��J#�����t>K=����A�K��u��ڥH��ɋc�7	F�̑�7�����ܯ���|E-v��lH�q'���-6l"�z�O�cc|��
�� ����PfR%	��:�ƥq�vFY/%�)�m ���QZo{cI�q�!�"�χJw��_�iv��(��곈B�0-~Q�� �)��	U�3��A�מ`Q�$��� �o����љg��)X&J��8?��c��p�ҌF/�7�Q逳�f�쏼�8�)�J��9�h�&���@a`���NN~X��t��#�V��\�~j
C����f&�����}�G�Zj�~e�e��;�X`�T�!�z{�JO��]��k�l+�}�$���y��|�i�~��Tw?j���tgS��З�g#�%�'Fk�C�c,��qG�o-bH3�%nː���T���q�J&�w�#bx�w� �3�����r���$b-��c/T9?(k��"o�~�$�O�o�ܱ²-筹J��X�t+�2ɳ'W8`�r�-˝��G�h��A����������qV��%��.p+�i��B���,\>s�f��=��Ctȕ����몃dd�����}�
s)R���Ӏ��D|���)�{+R���ʢ�2�债�p���;��f��?���컋@S�?�f�l,l8%@�n�8��Ze�� 7BH$`�t��\Q�X��ƈPK�@R�'^�y�Λ��h���װ�ֻ�ֽĀ�9��f�%�,f`凳nf\՝ ���A'��D *V�t�`�ZO�Lrfj&<�Ѽ��&��b�*M�c�u�N�nZ�~��A��j�]��h��\ ��YÌ.��A�0tw�߁�!����$C�ET(JY�PQ\&�r��lku4,�Ve�PJ�JpΛ��(�R��	�X�h���G��օ~<Eg��fo\��Loѐ���!��r��Y][v���c-~{��R(N�9�B�\�+�E�oR�#c9<e�r��f� �K�'.ľ�\'���1Vo	�l�C9�j�)�S`TT0�O��LsP�떞 B8k�Uv���[fo��ԕk(��vD�R��4���]$�CM�z/8�Z� �AVORn�
tD�����{fJ�/acN�+K�,���n�x�a_�}�E���3¾�d�U�1j��Yp�W`��;1���;�5�e�`�g�-��/��"·�b��)D�V�>�I�3��'��}���o�ҫ�C5��I�<�$���D�!�z�<Cγ���9"��~�)�Ä�z��_#�� ��2f����2�ek1�� ���NTb'ÃQ�n���?���}�+�������f�~R�?�7O��>C�ȳ�$deJ~�UL�� �A�Y�vb�c�����>�sJM�S;Q���3��Gt��(K9�����"r�*���G{��-���Zw�� ;j!���O�Q򪙖K|����<�X�?��m���Ɔ�mVZ���Q5����0�a"�A\���|76��$	���g�(�qvܑ ��FϙԶ�mW����w�[���:�ᮼ/�ra\��D��2��n�c$����9���8�q#F��)�
S&;�H?�3�G�C����0��L��z��_x�b���O�	���'�͟��kKE	�N+b�c[�.!�ե��i�I����L$����H͊*�\u�b�|doݦ7?/�43o��k��V:����KF�i���iQ�{��X���j���¾A��cd0:���M�.����}q[2��\L�|G$<0hѠXV¹��M���hPl���E��7�4��q��Ui([;�}��A v=VƏ��?�7S{��6R2a�<��P��.Z=Ա��YmI���)��d; �c�Ln�O����b��u�$��A� �q &��h��=ooL���(UP�_mRU���b�EC��_C��g~hq��y���
�Z�f-�	0e�t�,�޺��S	GT�!��o�w9$	�bb�{��Ҳ�Q�n|�kM�>m��m	�ˎ[���i�w�°�h�:�o7k32Ny*ҕ95ܴ��U�XkO�Ô�t���8�/�'�	�M{��8'��Uv�<��@Z���JC��'�s��֮ч�rm_Kߖ�'@�����l%s�W� �� 9��n�(J^�9����e��ݠ%H#�&�weS�`G�*�8�o���)�����*��6Ph�!�����E�!Ozܨ>ñ�Y[�w��31���>U���$�)h�d/��핰p�RLFS=@u�*�p���L�,CX���}�� ��
�I�lC��	�H0b5�����%�̟[�2�[�����t�u��y��������Q��g��:TK��.��H�X��l#�Ab0mr� ��i���2�KI�W�=�F̾�)���?%n��G��&����+8R:aA��Ų=K�S>�=Kg�pb0���J$�����yql�P��X494Yc�B���t��#�LM�b}�ٺ�$Va��V���ł9��Y��Iꣳ( ͡�a�����1���U�ы��/���ֲ[LX$�ک����Ͼ�!��-@""�1��	D�KoRcg�QY�{�$}�d{1-�>��ִ&a����}�踮L��`�<)C�S�pz�[|6�`?��lT|&a헖@�ul�Κ�KX�+�P�m���$x�v���PHOV�	�V�K���L�������ށ"a��)t�3Ly�},�2])נ�2�̴�\�g�?'�8"-Q�,\P){���p\����f��,�bmZp�1�O��T��}>��C2F�T5�"�{�o��x?#�<�c9?�;���o��e�t��m�u����xְk�3?�2G;C@P{{Th�$,P#���0�$Ag$T�(�Y�pq%�w��O�n������S�4T-%-���P���-� 9lX3��0�����3i'J��<31kR�ݓA�~��5����Y�^W�ҕ���4�R5ju��t
�92G����l��,b?C �U��D�[�L�?+�F���NCm�btSD��I�d�'���f8��d0X��ՠ�Y#A�_�]c���i�Dp�)\���%ZIpw�wy\`lt�+c�ɯ}3Ub�W�¥.�L|
�']�^�%��HjbY��j!���1(ʀgY���:Q�2�qva<��y�S����1.��)�T�I���,g�IeٚM����^nV�~����9����:w�-�8��ZBH��K�d����o]���s1(��U��k�X��I��h�I�ʋ��5J�όU�Ӌ��}�ڟ�\p���9��HJ�㚁�d̀E%��;��}Mdl�^���WS���τ�z�A�5`a�_�(ǳ�`)�r��G}R����B�K9� ��̈mI����I��.MD����_8]3gg��ԓW��T�#����7I,��ck�]@�jNm�r#���0����/�'�X��.� ���ћ �n/������E[�jԀ��p�U�o�ni�L�j�Z�� @��x�I{��~n�$�f��#Y�n+�##�:T~�^nT���Y�	�d+7�*��(���m��aV�z~1{���{K�ҧ�tîBDs��A���7��)��km�� ��7���&Z{�KЯ2 �"�=�@+���_��.���2ׂ*(b~�G����4�S"�$����.�Kȣ����&z0�E+U=�"g�/3u���q@t�w
��̅���kc�ut�T/��ݍ�p	��=���[Š�_�yL�˫7�Wk��!�ǁn���m�ʱq�� T����W=^�O�]���WՍ6.hhؽ�3���0�'
?>���;w�A툔���b�	��Tp���藄�����P�fHݵ��_��W����)�U�gzu���1�Hb�t֕c�����f7ٖ�(�Qw�6��qe�^����S�.y-6�ib��l�vB4�s `زr:�V�t�U�(���>�3I����P�{����2Hu*(��'n��j��%�g"�R�Ql7�h���;V��rF��ޟ|��k�U�~����t��.���n4a"�^�������MM���
�eEO��S�5S��խ�<�#+[d��w٘|y�y�����=�1Z��zA��B�L���:
�D���=Eu��Qs�Y�xt7�ĩ�+�@qb8�:�܇hv�M��t��ҵ��`�.{���+:���:�"ׅ�QPM�$��[����lG�����Çɟ�y��N�f��Ai�{����T�����29a�|K�!&a���<���-���N���r�Y-5׆� jQ=�蠣�5r�R�/�g���p��x�z�� �@�J�l��P�b<n��lXC<�.<���:�NkhUcP�On����4�����Z@̏��ؤ̮���D��K��	,2k*��Ɏf�_3u��u��.f�nߞ_�Xrlѡ�}��p@���f�6��3r�r�������,S6��r�FѾ~U���/�F�I��h�P�&$���9�t� ��}ܵQ.��-6���C�½�k��'�'�ͤ�r�"�
��{baeB`Շ�->�*�z�^[�a���h�؂���d��*�KAb+ܝ�i�������D<�;ǆc���({.�XD"~�����J�����6��IQS
h^�A�C􆳓%K�?���7�+>ƪm[��e?I���h��֔D4K+U�UM�x`.b	D�����N$��zk��B��,�VV�����t���߈�i��?�`����V��޴+��y�,ҙ��,������̞��\�{����[9��6�>h�u)8
v}&�G�"h�X��dh_���2r��(ϥ�*}��~�-6�\��_�1�t�T���<M�D7C=s-ݨGdq��?}�9��p9���>T��t���V�@+���NV���qbc��q��H�Cv���)��kpw�o;�"�)'a�$���k�kMI��3��Q�M������%�n�K����o(�>j�R��3�|��Y�9:R�Z�\��=�E��.��rDIU��̑�4�ZX�j-�eӎ�~�\��ī`�3�^;����s���xT�l^��T�-S"	�=>��0�b(�O�^X��f�#�V��"�	���v0�b�C!1��5����1���V*#wP�4�PdfJ�SR:7oDL��� �A�m��.)��Ǜ	��^��pQ~W�@�Y��(��º�#bc�4���_�8W�]�=�؋��i�,���K�6�s���is��Q�,)���UB���'�3_E��Lw�9	e��F���.0��bN�	O�~ow�k�C9�x�}h�J	W͐��tB���m�)��_�q��f�PI�΁�=�S|ߦ�r6W��FYm������?�pێ,�?@�~j Yģq.�*�,$���e<�p��$qf��o�ٻ�xEIoWO��x�,���?r�q�������լ:����ч"1�C���u;���@O�Za;���Q6�+`�n|9�{}gc:$�aZQ^��SF��V��5G�� ��5��is��K]PDqȟ�:0vѝY@H>����b�KJ�7��D=e��O�e-��":ݐ5I�p�[�4F�ŉ\�?^�����15�,K�@)|����������<%�mJ(�E\�شL����n��Ҡ��=Í߅���[c�	e9n��q��1o%��U>y�$R. ��|����Q��i)��f��?����]��Pv��J�y�MQq(�G$h#�4�)�+=�v�����c�$�$J�_�.�V	��t�jv}52QD�zʥբ��'%Lk�юb�꯬.Ά㍇�˧��:��U#L����r�g�OH�;�0���4l�7J���q�a=�c�`H�E�� p�2V�1�e����Jg���`���l)N�ԫ`����X�O,�ϟ��S����&+�;��ސEB���V<ؽm;��jv�v�˞�����MD��w��lx�y�s�
9����nu3R���Cӷ*\��"�[c-�;��yZ��w��+�l�>��`v�X����k�˞�<�7#�|��ͼQg�-�-:�5��cH�@��_�C¡F�jN�&��@�O�����쟋 kIN�Ǳ-�\"�:-�py����|�LM������K0`C�����֔��1��FB�/�.��^��/%Hfq����A�u���C�o1�9�����r}F5t����ؒgf��|C*?��hQ����q��R�u���7�
�!K��`h��[��v
��j9�D%?Є:�*;�L����)P+�1�Tn�$����+�K����u�i�d:�y]i%)���2���a���	VYl�v{=,�b�ݢ�����9LA��?�m$�kv@z���_�k*#�w�9�_^:��7�*�����x3�I�Q���Zm��	�p8���_�7@O}�YSxmm�J�6�^��V��������Z��]��ҜW�q>��s3���2|��??���X��gL"�#�O�A��6}N�j�f��5�C�	��Bb�:�����v��/z���l��?
��D��e��ʶ���?F��0LC�_E�8j���&�gd5*��R��a��W'�f���c��Q����Z���-h���r� bfYtv����v(�믧6�)���W�5\�{�M��ķþ��=���5*��$L;����A�W��h��XNd{�a�9�Ӛ�Bχ�U�7��kq����}C" �$�D��C|��9g��ImW��X�۽S1��u�Uh�+f6��ę`ϕ�����Yl�����bI���.���q��9H��.�D��l\���S:�ܿ0�j.O��,�ێ��#�C	���1����H8�+���QKib8����v��xB^��� ��|��p�	�IISb�G1���� ��U��}*I�ɯ�Q���'�L�h����d��n�g����r	>XI�����,m���!:)ս�D�`�n�6x"�׃�e��c�͗�L�����Ȕ��%��s�}��{��v��}@�%W�c�y�4����}�6��+l�E3�/pMa�X��'�x"�O�z����Z(YN�8���]Ԧ#����Hɱ2��H�`�H>x��u̒�uV�Q,���9��.P�s���
����(n�q���D%1F�&�K�@e��]�<��9�v#_E9�	��r�����=�,$�4&��s�KHӂ��@���>���Y�z�ɀ%�R݌����޸�;��!��!pg`���ٶ"��e#�>��/�kӣ���=5T�4��1u�`{�(�Yfq�|�����lm��K���i��F�t"�s���ݺ_{6)�u"�H1��e�j�h�0��s~�%�oK��X �~/+�m��½�c[��p�JD�R���&K8\��%v-b���Hŕb��m�|/������������tV�a�K^�&!.�+� �Ӯ�㙖L;p�<N�m�䠏(x�T���_��M��&q�z�i�����(]�W�<7�v���')�x�	��z���'����:��Y7���|���]K�ݹ�ߊ8_;y���gNo����+����4O����%�r�'�����r4\�-�
�%�O0UA�K��N4��X����D��t�b����qG�u�W�</��VsS�-�j�W;Y�a]�ED���5{W`�'�^�(��"ɺ?���ܪ��9����4����eh9ξ	Y:�k΍i�z�h�0��%���<W>6����Am��K��>H�rq��lt���L��	zͲ�٨{��$�>]��n�/F��a30���krX�h���8������U7I����Av�$���E7~�^g��>��ښ�< E�>n�ƅ�'É�̈�������d�h��,�ǰ�R�,�Ͷ�ت�&���ąۓ��[?�^X��J�K�~��W΃>�K��� ��p]�x�����4G.$ kPY�����Bj�ݮ���D�v�7L�"����BR+~��sn����*�c��8��O܄_GK}{��x6:^|�]J�������+]J�ΎI�������&!��MuѼ�N�j��Ǩ5x�"p��ۑ3�g��0I����Uk�t�O��̢C]�L����H݃Q-��4�_�?���Q*�5���r�-) h}����M(C[�M��'����:��UD�FZ�v�3P	��x������}i��%1թ/;���ܽ���`��ȗ�?shn#]G_t-Uz:̲����*$��7J2��I2���$/�����K�h)s��.&�0y�f��s4[��s=�w�����WQP~�o��Ay��BK���=O�A���~YC5u�&��g�)�C��Z�'6�Ox�������� �B�Pr?"prxQ+W-%y��$S��/�C9͊%iy��%�):K��y�ʹ���C�O�
��9wW׹�7:�+��kX������3)�A�����N�a0Q��+O����~�Bo�<k؎���-��ׇ4t�)���{L9��Qq{�
���{����Z1_�pS,�X�~Z�&K��!_���EqM��w;�)p���S�|��w֜(*f�sp��;��(��}��$�"��/N���|��6�g�=�6���'����dl�'���U�=%�wQ$r ��?דh4L`$��V�J/-�:�!����u�T�o�|�cm�~��vܪs�1Z�0��%�@W��8���^>^�qh���ޢ��Jӵ�-��IN�^Kce�5F��?�5.��q�rd3&���Z\g����29
�Δ_��1!S>A�#N�x�oӉL�#�2���N͞�����D6��Y�7�K����������<�'�P�Nto���$��uY��b�H�L�&�>�Å+����Z �����|"���y
��ōel��y+�����Zo!<d��ޟ�ζ�2�:��Mf�F�
�n�_��(�֨����g���}	��(7�FpS�a����C`BpKB	��b+�
ŋձi����V�4��蠨�˰��k�g�Z_�ej�e��e�Hwo��hq \*�s	�a@�3.��s#cTD�����b��Jx���U7;��`�MD��Y}Y�:l���w��b���]���I�aާ���@�Xm��F��ͯ��Jj���7UXU+,8(�Z1����'UP70�
�r|x@�Z�>�n$e_��vE�$��������w��ଆl�P��K�\��2Re2��`:p[Vhn�v��t�=�����J�YP�/�hS"5��C�ǯ�A��.�r�ҲY�>+:b2N/s�mw�]�?9İD�HI��·�峼#2N�2���TŎI$V,�A��=y���YZ_kV�W����uP	��.�e��Y�ـ�4�Dz�L����P�<���؏�9 ๵�ݜ�k�8��E��l�պW��G�G`'(���c�:WrC�|"������z�m��s�����@�2��غ�Z���vc�F��[� �j�S�S<��d|T�5ƴ+�Q�1�OW�
�^e�6�P���}���y���|������!���H5=���6L,�@+�<�I���e:�����-�b��= o�����	~_���E��#�G�z�gp��b���B͓��m�湵��B�����}�&�u�2I�`.7)5�[��S:)�a�{�g4��+&�$y����p+K���5����1lg^���g?����!"��	͚�������vĥl�����E��Ц�D�Xw�B�i���b�FţW:s(���;|c�Zr��.ɻ�`�6"7@#�>������쨘{�=4a-t�_4B�˧��Ƒ'�䕑<8S�W`"j����xP��0�����V�V�u�4M,d�G;D�M�
x�"��:�1������W ���*|�x>~P�o=��Ȇ���̣T�z��2o��7�r��6T��+s"��LF�/"`�E��7X�x�bk�`zߒ���
�wWQ���[�4���\5�c~�@=d`l9��*S}qk�^�ߤ0Q ��-G�p24�	��#��(2"�ܦ��L*��cl��ǣ��5�9�O����]FB�� �l�,��Iθ��^��aڃ��-V?8ZY5)�X9���;�R*z���`ݘ	v�����>M]D��O��~r��I�NE���~;��M�����[��$Zt׫����&�+D�""ռ�u�Nc���9��n��֋�(���9���hhJC �����|����u�/`LbE�\}  ��k��	0��2K��
���J�\����ηC�vę��@�i �8Eņ/BiLK,ІK�>}�و����&`V7_�T��]�
�O��m���b�cD!�� 9N�8BkN�-���<��}A�L|9��:�Ė堘��L�a���i�����ֈ��MA�<�/g�K��Zt�3X��LUeu^DH�
�a��sȋ�^�U��{����7��nAǽ+�m= ���g��fU��|:�]�5f�m5���������^<Y���ΐM$�ac\��̟�rr��U��g���3��:(��Ř�i���- ���N����s"��*7��u�j�{]��CWA.���'|�m*�H��\�ȋT�/�+>�0��`I�5T��/K��n��V�z�o�v��Ud�w*�Q�&4���㺷���� ,xS���ݼ�m��G8f�ߏأH���Yh�36�($8�)w�^��H �`��RL��v�,_��z�b�XƊQ
5A�'n��_�_��t�YCb�ʱ�M)����q��u���F��?j*%��[]��-bv�!cλ���Gc�)�-�hr.v>���B3�v#��ژ=n2���,�_��U�73�i��yq
��hA\��lC�L��U�uݏ?c��D�1S�53F���->7ѩk���^��2�
BD�T��������*����z	M*M����?ҍx6�<�_md��&!-�&�mEY����u�g�mz.�2m����N�%�������9�_ҕZZ���V;#$�6m�����uH��β�3 nI}�,��2d+]ir2��4�gD�T���d%�b$�g[�u���A&TI,3I�>�to�h�ږ�h����Tk��|��.	�x.�tIl�8�&����o���.��to�Y���r���� L*{�[ࡸe�N���n?)V �a����w����#����l��R�Z���1�в&�aϡ[��/X�|=��z+�	;;��C�I��4n�-��;�nDZ���_�.�̅�&����HDl�'���-����)Xc&����g���h�=��<�Y^�!�p�ꈋ�K��G����E�����q�v��0r'#�������[��FI�AݥzI�������@y7%���|;C�a3_��-ܳW�9c��|�$q���?=8���Y��_ׇ��a�/)��)Ė\��H;��E�Ҍ�H���x*��0�%��K��{�6q�|BM������o�c˻G�h������5s�x���!�9��I����Y�E���
�n
`�p��+�[RJN1����K��Ҭ�y���gԷg��=7�ʚ'!�q>��%�̏\��H���R� }�a�E�^w�:��:(c*,
�vG	�`Gh��4�녷 `i#��Ya��?�k4qD���QV戒���u�ߛ���� h��!�ǝ��H�0o
�(d�_	�3��#��$9(�h�J@Rfq�k�=�Bo�l P�Evyf��=��iKTƉZ�.I�E�6|�#(V�ٍ�nef��":����C�w@Qfx���P��e���^!����Cq �mU#�TR���2Ku1��a S�к�B������x���隄���=����������tH/�����k(�5�'�0������b��ĦN^�_d�j�[��7���*�?�I����H�>7��t���^�����$�=6��q�g�q-�1��6h��6c�(�.�9)�ϣ[g�v+/�zK�\�/v��Ď��n��6��EJ�ګ*����lGŒy�ik����y>�j�yE�;�l<�տ�;���br�<�+^}�X�"����a�e�K�դ�1"V]Ƚ|�P]��X�r����g��������'dH�"�R���U������������%�w:f�W޾�,p^x��� �����4��^��p���+� t:0mε��!�6���n�[R��E�#螎�l5LQ׃|�V�&\e�ad�aB޺t*��ˉD? ��"��~�($c�J҈�^`
?���ǁ�����G��'�u'�$#~T��7�?\(��Ya��̖�m?���k��^�*Fb�G�<���.�\��9��+�
9T�mhW?��vO�K�D"�3+�f��v�����~����ي̝z������ԤX����K	�d��Q�F~m(SQ'[L_ۑg�<������,U{��0�$4����v��Q wU�bGW�\��6��P� ��L��^���i�~UR?:��{�����X�]����=?6�Q�}�GW��Gc���"h���k�n��j�Q�P*Y��J%�W�h�	��t��bɹ��W ��*�Wy���/�4��ʄ�'���ކP�����L���<rp;�;�g_��B^m�=�wڊ1�2O�V0�d]��{���\զ�ϒ	͘.���d�Ҹ�v��]�{����kD����zr�����Z*	��A�X��[��2%��eD�c����&b��2R����V��	�r�H2���#��t��V�c�w,��A?aO�n�uN(��?�
?��j�:�7��~g~ߥ�o.������[�y JHc*^Z�0FG��W.{�P��Ue�϶�P5dm�o! ��4�`�����@#�z���+4�}d<C�S����Ζ�P�$����SZ��>]2dD�tS�&Y�>Z\:�	y�D�4)L�\SP���Hsk�s�C�36:s�|F�>TjL�U�%1^! ST-������T�+l}T�F��Bb�r��V��my���W��Ý�m���\���!]����������L�~�ذ�i7���b��~��xg�(�V�{�bh�O�#�����1�����S��"�(�8��;��$��H'٣�i����p�=���M�ֶ6��Θ[�B6����ML66RUΝ嬖m��+�Xv
�6��\\���j-;��1kZG���2���)��˔�X�ն���A��"�Ǌ�F�����?%���s��3�ஊ�������H�1K�c��3}2'�rL��}N��ܔ��?�?�k�m��
<YgU�w?/e�xߵ��<�b'a&ϼ��Wd��F�%��j��+���4Z��ڴ���{;�x��==��\5&a2����kv��˞2��$�-�T����*O������	��[O� RE�!��b����%�RLQ�NG�(�����d����{�n�%/>������Ƙ5�܏�ϴ��3����w�?�p�=}�&Q���-��w�����3����k��LҞ���%?�ӌ+FgVX1b=�5� g�\YG�0�k��8���;�1�[�iZfm#k.���ó�~E�+���e��x.��2G����hݻ�vگ�(�Q��T�FHMز�V��v��J~��DZ��X�Y�3�B~���"t����2�NT���Y���
C��N�O�?�Y��������S�4�w�K�K�x�ԯwN\��ʇLXu��ŝQS��ML��K�u��O�.�{�1�w����1;��y�/��w�g����7�[��'.wO���5H~K���x��&&��iGTݶ?0����8�S��Š��Sg�oW�����T��@�9������T�ȯ��+���|�	6lw�m�j��9������C�d�y]�:'��h8��j�;&���=�0�jٓ�ҥv���.�XCw�@�[��!��-J�#CHh�r�|�C�
=�Xʺf���ِMy�U�R���2zҾ/�	������z��}��oS��ّ�9g��k�hqx;Ϸ��R=�_�o��/�鴂U���Qa�Դk��R�lj��9�]	��R8��-!ͿF������qB���ؗ���Y�N}�R-�����������|�1�1"g6lB���	)쌼�"����+rpL[�K0y��i���&�- ���\7��j}�����vth�z-�[��pњ~���X��K�d�`-lC�g �&wD}���rTwN�9����N#�7a�"t�F��H����E6[އ�OX]���i��3����Y�ћ�B�UQ[���r{�p�}N�gT�*��R1=��,L���@����� A�u?���n.�9,��n.X/zvH�����+͗�w���(8�{�5 ֋�ǏZg�/�_��+9d�X�)0��J.�U���K���WVje'6P���N�������,���D�I�p�X �(���&�[���҉�ǅ���/�'&N����|0tB�p�=��-��\_�s�5V��[ճ��&l;���`��Ω�Ն�\�\��1�q�H�{�g�3�4@������//�E��/��D�cD�$�59�$�&�H�k2As�Ze��:���z��[�D�w&����x�Y� 3���B�;[^C�|�u R����9GE��~d�<˛�Q��0m'�(���o)@��7�;TЛ9�8�r%��#ر���JU�#m��Lm�U����al����j�t�c������&,=����'@X*]��Y�� f���I��<�~��m �u�`�H�"Cw�_x~�d�A�e�g?�7��L��Ѻ�1��g�~�l��h���m/���)��܊&_]d��K;�9y����M�(�JD������jឰBz�]qtJ��gJ���n�V߆ձ3.?]Q*�s}�;�q+
��	^$=q U}�6���VOB���l8a�E�.��q({�����jG&�N�̞�S�T�o6�����[��o#��W�q2�>d�H b���DY�)b��(��'>��g��j�����_�Z�8&���ky��$��� %�kJ�����F`!&��)��O����H\�>ܙ�:!.�s�[/lڅo�IP .����K[����%������+	9�.T3T��7��mN_���_�E$����u���;Њr����s���O|�����n=��