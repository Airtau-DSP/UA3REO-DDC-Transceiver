
module debug1 (
	probe);	

	input	[15:0]	probe;
endmodule
