��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O�u<�9�F�|܇�?g��>v�P],	���J��Ӟ��Op[�Z�rSCS��46d2��B����ȩ�� pI���Dx���
(�8N� �1E�>��"�,�)}0#��b�g]Ƥ�Z�cͥ�5�#��ᡑ\&
�YH��9]����-b�N���=ɟ��t�2f�Y���ۉk{�x���@՚��@u�-k�Ʈ�[H�A���B�QW��ad:!t70�9HK���װ��;F=��I���@u*w��c�.�c� _�Qջm	�/����J�A���͗}i�/�V���<	�����c�=
Ц�㍊mSY�׏�� vU�ߍl�2� !F{�(��L�V�6�o���Dz�z��Z��5&�P<��a�4lp{DO��s�:�F�搿Ob��ȟ8v�$�n�x�J��^}L�F�e���b��h�����. �$��e��0�����1�	�ir�=�ɭA�JL��r>�#[�W�@�jv�k@y�ەM�T|un � �I23��f�I���=�h���{��I���B��?_6�b��.%���I��׹���ѿ$g��F� 8�����sU��D�?�d�R���կJ�69�7U:�q���S��bk|�!�-�(,{����d_�#H5K�A��SqI� ����6($���2��lrϷ��mbB��o &�u��v��:�hn	q�^�Ѭ��q��s�JW��&�	#H�K=q joC:k]���8ګau�|\��w��v�Y����E�����N��#��O�818s�)��&btk�-&ge��%:Z��A�B0r䜴��OI��Y��s�ɛ���'��6CxB�`8r���C*��}��������(��R;z�(^B1�#M�H�>Jdf�j������̢]15���*����Wdj��;���I
�͵��]�\�_o>�6ĩc��b����G�&+�����c����F�,��"{M�>�p���H���SdϢ��!w��nHw���c��ccs�Hi�8˶`RG����h������,�S��PX:���h���\
T�8�(M�ә��i㽞snb&Ya�t����G�簂�.������!����� z*D�F�@�Pq�W�m��3�<���Ğ?������