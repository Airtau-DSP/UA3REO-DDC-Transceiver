
module DEBUG_ADC (
	probe);	

	input	[11:0]	probe;
endmodule
