
module DEBUG (
	probe);	

	input	[15:0]	probe;
endmodule
