��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k*(\&��Y���z��;����1~;ó�!E7+ Uߟ �v��M�a�v���]�P9�Hq��;��p3u*���)a����9�w��mY(���Fu���u8G\��:��^��_eb��.ڄ�f��h��(J���?�G����-��vP���y��+c�Y�����=q��%�h*���h�Z^��=3���f����8��@@ޕ��`́�޻��=7*�K��vn�餤6��
�}�����L�ۯ���fZD@��G+>�=��V>?_	��%%Ƿ�H���6<X� }��f��K&v0�otE;nP
<�:pf:����Fp�p��[�<~x��,�&�z�v]*�UW���~:�Z���r·�H 6�h�%��0��!� �;7�!��B=�JX�G�����Af{\�ϟ:z�}�(u�����2�;r_�=��.�;�5�'�)�p;$�!�@�G��)V<)�����g���ʯL1]:�Qm5+��Cod�����X�I��ֻV|�S¦��ڮ����R3���9����,m�M�E]�uf�?@��ɖg<�U���U��,���һ%5:1:��3�AL�ּ�w��DM��o�6`�d�L��4а3	� \��Q�l���z�����}#L#T���e1��4h;��pǠ*�����H�հƤC�i!ݣ��ݵqbX��{�'j���r}��O�w[R����kB��~�>[#T8��ڭ�y0�ߎ?��p��H]YO��A��M��B�n�iz�[(��'�ve�s�n�F���V��I�2�?Vw׾z3761F�h��8�MN��k��X��~��[�pH
t��rl�;Bs$�q��s�z��:}��	��D����#�7G���f���
�G��;�����/85��/ ��ɰ��y�|��5�����{	bm��AV��g�=�ԁꊕR3$��n��L�wf�w�!믛H�!o�=j�f�$%hA��gn���s�������9�?C��U���5L�A\�7�����r�F�c���=$�C��:���zZY%���qO�6ՉC��9űY)4k�|Gp�5�馓AMn/O"ㅔ��C����� ��x�����4C�|͊�m ��#�6e���o������&m�p��饂1��=&��]����^���@��_;!5TԽA���֜�oS#�$!��*��Ԕ�RX�em��ky���,9�`9ʰ��;K�C|%�d%Q�'�D���4}ndaBN^Ʊ����V���m��[��/[���=C5%5�HXȓ��^"wetN��8��#	�����g[�pNY���+�Up~W+���rZn���kw1� ��W�&��~�s��0�O�vj~{%�>��H�=�s0^\�X�H)��� wוM��E���М��bu���(�Gގ��$�93�!>�"8!Z�erܩ�e]�	1���R�-F;���������-q��혓����Ocw��Ĥ�D"=����{�4/9�z�x��(���y꺻̤?�,kDV�%�㮊5#�&� O%�k�\�X�#@�{�����Ȳ�:�cI���1'�%eջ�뚻N0�zO�#��V�\�.�+�NU���N,_�7�sR����;0�f��'�D�(n�J�#qí���V��]\��z���!�	o_��q󲝝���J���&���q�Ͷ$>��L|T�`�pD���	��!��|��������;�>/���e֡��R?�MiY�.^4�:jΚ���F��:&.���!�me�LAS��Q��S��ĳ��b�|���ϱ��D^g]W?H�Q3<��5	3�#m��>�y��*5\�BO5�Ί+�PG(�I��Y&G�D(�}ݢ���![B�{�B��V��&�\.PH��W$����^��/��r�ˆ�q��HxY1��b)�<ey���R�S��4���[`h]�n`�E���+�����?�k.���iYK�=m�������o���p�MF����Y��0�:��繽\�;�g ����]*�ֆ��I�U"���|3�����
�]�*)� 2t��@ ��M���B��)�h'��̍w�.�!fP���@�R狎c����޻�7�	l����"�<qO�(���w��a���G0'�1E!�F�����:p���`�����%S�q�<�u5�D�c���l��AD�4$�����ʋ������I��لiH���,U�؂�cE��PV��Bɿ��2K,ƹh�pGVe��נ������}���,�$�h"��8b������t������?>��ܟ�5$���"�L�Dv^"� �#酋!��2'�!Ȩ;.x�0��P{�����1���qBC������z��
�!u֛"/���A�����d�i_�WgS�+W�����K.(=3<S� _5���K�Mp�����Q�o�t�M�����r�~-��Q�vɮ�q㝠�>=�Gń2%OŮC�HZϬ|>H+���V@�_վn!K8�XGD�`E��|�@�F��=$�mz���'�4�йn�=tρ��=@"9��
�-&*�#T� A�J������,	���\�9ʴ�ah��n��+O�Kp ��Ϛ�+$��j>�S�t�d�@䫨̮��-fr`��뢞��P���3�<�&�x��l.
S��Ě&sc��Ll夀A?w�U�r�d�c�<�+xHh�v�������K��0<���J�>�u�(�Ga�W�|߲W�aWxc�]�c��|R��44��RP4�q���Q{�&Q (�+=��Ύ�-!�Ao�[�-�I�ǎ�X�V�D��kIӞ)�����4ϸ�������܄a�_X�Z�GӠM
 ��I�)�g{�TNHˇ G�� S�(qs�n;N�CމU͋�d��V�����mޮ���_�jڟ��2]��C�,*chJ_et�KaroaR�t�8s�0������r��r��S���3��Rڲ�[�e��9���ʺ�����V�.�4��m|����\6a܎�|��״�Ԕ�v�$��_T�vckQLz�m���_i�XW��d���Qs�!{!���2���-�Vx�A������p�5���Q2���O�4}��!2��W��_�(k���'j[�X3ȥ˰@?��g�bGs:��Z��������nB�T���8ýA�n;�^zc`���-
�D=P	��nĻD�p[; =w�eRi�S���Z#[/���e�5���!�)q�lL�c7fH��{�)�Lfܽ	��v�����8����54q�_�I�f*��}p�|�'�1���ȿ ���E�sq�XH�C��ܰ�)�E�⺼Y�+���u]����'�r1�3Kz˫����q�X;�6[f}{Ա+��-F��Y�	P�D)0�	G�
tK�HT_�#@�Kv���朱&b�|�-K��?r�2}2�V��O��&=fl�H��g7�E��̋�o��v��J͗��xL9�y L=�~��^���cՂ��w~�V�96�O��zs�2 �m��s�y��<��ZsS또5���?��T.���_��/�Ѩ�\�������LUn|��N_{�D�gjU����Sg$��=�E�seg+#����m�J;I̋���ݝ#�ޔ K��6&�'ء^S_�v�-�Xp��e�Y-+��'#�k��������+Q��T�w��u��ϧ������J�B��'��R�NW�xP2��b�T;w�z�ƸI�	��a�����&��ޗ����﵋�^=AT'4&�!��,���K]Ն�����+-%�+�>�9RN=�4����~�ۨ֐�0��0%��r^2�=
�`*���죱d��`�$��w�zV�i��E���=��;lF�O.��jH�k3�v;9P�1{}���,\��-�>)''<j��5�^�c�G~����Be���=GG�+��	�h��OH�0�+���z��^l�rXX[�&�R���O�a���Z����}dI@|aw��7�Hr�t��J��$񹤛���&DC��	j	G��K���&�(�9��ZXc�g~�\�� t�����a%6}mok��K�����a��/������E��dI�����a/�Y����+��0l�ppm���Y�s=�'�C�\,-~��u���i��*�M��پ��EMX*�]K����5"�i���]��6F���զ�K��g4t��ы�����ժf���0%��JE�*P7����v~FH��R�j��e8!��i!��-�3��ؠdAP�|��5�U�w%2�b����x��Nu�f�tր%H�=o2Bv�| ?�/VD+T�E`x����h7"U!U�և����Sﻀ�x��b��Y_XF��	OO"�M�
3A�_8��<���d5�c�@�`�� ��D�h*�T����|���ϛnǙ��-��~uM��x�����S�j�sFB�X>�7D�0Z������tRe;R'C �!.�%��D�w^D�k.K3>+�ū��!�zC�.2uE*�0�l}�,{��(���(V�؍k�e)_�U��\b$�ܵ��8�~��X�_���Fq�‹�	R�k&��u�O�.B�>�M�Yk��0�9m�^h�:h�R�:8�x	���/��	!*�%o�(���ލ�1��qp��<��{I�S��8ӢE���2����{��`_fx�V��a�E�zM��I�2p`�7.2�\Xm%zg�2u°)��E�\Pȗ+��Fe�~��|VO�w����!9d1��ͭ�{�,nZ՞�յ�C�ﶂM^]�t��!_|�ީ()Fn�J��ݨ��r��O�1��1�iS���ҳ�bzL���7�/ni��.��ۏ���8\���j��$7Î��"wNn��������p�a�Z8�OI�)�	����$�����0�誆�Ӓtc��=�[���Cǿb3�*)*��ڎ7��v�uF�%J8��k�~&��v@���˲�:������>�7�\�������8~F^o�O��c�����8Z�:j���'S�zg8��"U�ν�J��  #	_�+�K���r�1e=�s��5�֨(�V1��9�����JnI�a��J=����b�ng�>�>���TKԁ[�f��J��o��3v`�]+~K��^�g�㢨ʅQ]����I�f2���T�B����ᬆC��VZMȁ���P+zLX$ߟ������D�������@r�E@0��D��0�xA=6�\�cAz���2G񃮸#�xL�y��bD��"�W�7�T�c�	�5^~�v��d�p�r��3{ʑ�@�K�]N>���	ݘ�Sj��﬎SA�a���w�1��c6�����mQ���0�<�PF��P��6�cf5��pIW�u	�*r�TLt��TS�+���as�+iJ�nV��ח�\]#��r��w���Lu�_�>#�B�|WL�\`Q�:5�Z�� {Di��w�hY�{>鄰Ԙ�!�Y������H��!�]��"�19a�K^�J��)����[�qVs>1�>��@�5G�+� 죗�@�KM��7&�@=���-b���'�R�# �*o�3馍��S 
�����Y�dC��?|�;��p�'���.��ت;��OLڞG[�"A0B�k�pE�3Mhvך�Gzn�,#�v�ϵ�K� ���@
<��.����G8�=b����-iW�LW�#XJ�+D�Yp	K���1�Z*�<p�:%�=Zr�<^�2ݨ��Sk�:e���Ӑ�M��r��/HL|U�2'�pakk�?4�l�%U�=�b����Yz��L�k�Q�=h�.�N��P?Xh��֥�ʓ��PvF���"�9^�~~=�D"W~���B
_TFT ���S4� ��c����GZZ���75(�<��G���?���J�Sx��� ���gLD�i0s�{�l��|.6��koG��<�>����@�΍���D���E4��+4%!~EQ��S�W?T)�ܑ�=��G��X^@��e�,����1E�08�`J�W�E�xq&k����Q�M����Q8��I��I�bIx#M�=�ɤ$�V�B�F�`yTCP20��uB�_@�n�l�����4+nD�C�K���>�E��a�%�(�^=o�d�(��f֪DSn�W�����JZ���j�� ��k��,�B�51$�9�{����G�ȕ�.���X�Qrk�==�2��F�5rὄ�;�Rs���!�