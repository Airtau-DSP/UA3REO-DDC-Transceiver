��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���'�ʞ�~|�A`�U���k�,�ܻ�zc����9z�n#�?Ff��w�Ϯ��^�����[�0�=3i̬�S��
5N���-)�[IN. �b5
��N��@<�"܄Q��X�q�E��?���^�Fǈ��������0�X,>�|�)�	j���%>�CaؿQ��vI���7�K��`��r��NA���x�2C�>Ɵ����ޓU4.'����v�X �n�+}ʚ7��o'��نr����]Ҋb0�����>�_��E#�C�W8n%nT:�W��Ҝ{汵�h"e��U���vd�$�3���쒘��鍝�5��SDJfގ��~�9��Q]�2\O!���SG�S�
���[��n�nR2�l`�PҾ����U�F��ӕd"�@�#4����w;���:�`�R�!EƜNn��
y�W��:�t{�/�u��764kWk�
�Dw�H?)t�����yF���x�Lh�^ѨT��2�aӣ�FÜ�@�&�av��,�'�i���� >˷1Xi�	\��) �?����ܕ(pT.�'��',r5���q<n�Tw 5���<f(��B`@���}CA�����zS���C�Lssk!e�����xG���c!�gb@���!��a3m�������E�fb�{����Vi4w@xh�/�82����z�Xw�kZ6�B�=�e���4�ӊ�T;/�|#���o�-OqN��XY�̢h��k��E��T�4f�"wAEQ����`���.�׶�ItM2�Ч=q�y01�\D�
�R�|�ߓ*�e#��������{�0 _��TO�W>�������,g-lo�6�� 1����d��M��fY�)�$�,�ߌ*N�!�H�)�򊰟�!��[/�
6-�(@,^@�-�2�7�2f����7��b��:�� �$gU���gz�aƃȣ`��LQ������K���y����-'���dNJ�6yaǳ�����q����ĭ�3D'�*"3eQ�M�H��e�����M��7>����3�ޚ�iD �&t~T� ��U�:Y߃����^��ǌ =���BV�n�`�vsъ'��	?$I(��A�3�Y�k�֪��x��8���Gj�5v.w�JR��(��EzXІ��`c�N���0��� N�w=ވ��T���n�3�;'���Yΰ\R"���d� LZ�nA8�Oj|���2*
�>�Ncȿ�H盍�� XK�V�j\����?����t�qGY�SPvz�ܫ֖�8Ϋ��=ǿ��f��q!�6Z3c_������V:�C#�#�vfq�ԐB��R��J!�}���n�����	���ݏ�=�&�<�ݔ�h�m�*��t�bfߺ��^+wQXͼfr�����]��$��i�%�7Of��;��J�_4�z9���r�ԅ��� �p/ؼ&8:gR8�r�q�����큪'3���;�`�E��*�6JM�� �H5��
/O���ѵ�8�J������= ;`���:`����/���3��� ��e<� r���M�-��Pu�H5*�b	��.�%ڦ���&S#o�� 	?u���x�mt��9�NO�=�� ��^��m��X���Mp��U�/O���������d��)����R'�%i�E=\��ק�<}�"K!�d%P|��zŚe6*|ER�-�F#���(9j�ٖ*��P~^.