��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����հ���y��C��wC������,�YՖ*�t��ޒ0�c�`�"b`�X�D� �� ƴ�������"����}�fV]�PJX�ુ�zpr_�BMÔI.�{D�,�,�W@���K%����e�㐁����i�a�	�]�ǇA�xO���٧f�����s&�q''����|\:�t�����O?��e���;�uݭaP�$�j����[�*/�y��:FP������h6�l,�VW��/��'v�g��w~�ל�M  ��H��r�W[b�D�|Z��o�N��qN���|t��<��?G1�F�/s�
��QIlP���P���;�Y1��i�+���C�.�7dڄ!gu*�7�M�:�^ܕ1�.;ȭO[<	��/�>�� 3P�Q��{����݃�ⓒS�џp|�{��l\�r�`�f�AV~�!�Σy��k|�?C����@؏:S�����c2VH�uɐ�ݓm��g^����Zf�ۏ@Ψ���a�}`W�N���Ӆ�0B�vзGܗ�~Ӣ�[����P�	!Z�������<ks���#�]C�;�ϧ������-��i�ZH�A�l�z[,��;L�2�rjo8�������d�M�2/��qe���Ԭ�p� 8�\D�k�@�[V��0��;�$<#��b�@0�.��K��g��(�P%ÜHNoc��N
��Ipݡb��6�l���!�}z�v��l3;��°sxPi���'T����WR�����`��D��ܐ�Ɔ
T�Xa_i}�=XA`Q�$�>MeѨ�isu�a�E��!ژ\�Vj��O����o����˟�W�q��PjO�Gf�k��M��Ǐ�h��VI����㪖�/>*4��B�|�*Od-�ly�˵�8����y���b���v�]�{]��> �?�]�j���?�%��5�
A�0�X:���\�ǘ�Bv�������&`6`�3�wh/�'+5ͩ�eR��iD���b|ME�tb�MU
��t���A�,��>��7��o� � ��lS(����Ԓ��zcT�(����[��f*��S=%�u���o��5� 9끙a� ����!���r���|�Ktm�P���2OĥH���Q�.�{o�_N8*��#�g��e-�i�#cqӮG����7�#�v"�|��Y�R�>�wݾ����m,Oi�,9�GoZc?^ջ��pXJ3�OU9U��\�-^ߛ��'�ʅ�C/����ϩ�}�Vkw��	@A��V�֭��,Ts	#��b�� ��HD�խB����  CWM_�����1�W'g%e�h����I"4b|��EX�:FMO��.0]f\ߕ�dl�v\��`]㦞�f����Z"�ŧ���!W6P'e�۱p��Ӈ`�r�A�+�n�E�r�B@�'n�����ͦ���5��l������ǸՅ�ˆ���<�봚�h����G ��+'d�i
��%�OΖ��$9�i���������G;{�f��+�����:���{ڐʥ�|��h���>��m8t�Srj*1�O�������� ?�A��U��o|�֥��I�$u�����ê��>ف�<��s}F���"�'6���; ��E<��+?K4�|`lX!�C�r����q��|M�&��k��!W��rD7�X�%��ub�+3W�
2�w�O�Mr�B_6pš����.��éZ�}T[(�d�;^��1�j<4�r�E|�u͆1e=}��G1�������[c¬Xýg[{R�ܑc�.�Ju(g�y��\;Y�a�a���{
��" h��Y�m�C�y�R�
$����F}�������	`oj��_N"�e�t����do	#H�̄;':i�L�@_�1�
�I'J��8 r�ef@��x����;�Y������`o�ɾ:˴p&>(	��u�)�8
��S�0��<�k���������!#:�$m+!�i�S��o�\{�J����(V��$ Q��3��*��CUo�Li�gt3��x��ȋ�Ɏ�tŻ
_�L�� �g>/���
"�+o���-CZ�Rк*���s�p8��A|��!Քd5~�L&7����]lq٥=
a�`&CUB�J��2�:�F�S&IHKA��&==Ku�-cG�[^������c ���g��~k�r;���3��x��ꩆ��R�x�$i���2L!��
�p4�>?Eᣝ��n��z|R7������=�lVC�`�{8���܅�����H�,����?s���7_������Hue�E�J�m������j{����F�BY�����Q�4o֞�[;hBȴoK�[]q^x�1rh+��}|�U�x�6��zDzdC�Eü�jĵ���IM�������4����4���Zi/��I�v�D+� D�`�|Ŧ�h}!5M������M'�"Z���7���Ԗ�ٿ�c�v$5�h���j`�#�DiT��ڐŐ�CwG,��k�Z�E��^4�].�J3+�T�����d?��/�kM,Wp@��oi	Z��qZ�cCvH�m� 6�ͭj��G��y�76�Ț��	)�:��1��j�z�R�����ڱ.�3��1�-j >����G -�bC:[�[���J��!Ǒ�B�(�/��L��r�I'X|���r�	�`��yw���މqh��r=�Ԧ��������u�%�0c�������*��T��^�*�+u���S�݁_��/��m9>�8_4���'C��=�� �<{Mf��|�\Co�t���%r�
�7�%3ǇkD?\�I�l�W��&�n5�X�ފ\������f�?���D��
����݄*�@�6&H�g@���[}��jd�����B^EY�{�no�َ>��d�l���B`0@U�⫨1�i����,P�O�+�$����9�5��H�s�A�fr���-��W�Ɇ��_��/	�灰*ײ��[���tP�/�@��Ӳ,m�kN����rg[sUO6�Z����d�6C-@~�ʷ<���se��x�BV^F�	r8��-��k��4塩!��,i{A�v�h����]*ڨoe8�3As�b���4��Ea
��_g+����\�7�1V���h��|��C�����e����2}��Y���+o߸��V�x����.bl?�$���Z�I���ui���c�jh�4�m������
K���&�Uq��.��45�x�pv����o����n|?�~I��T�p�1�V�ӕ�y�&qX�NmM��'�(ۅյx�|^9Mpǽ��(.C~Ԛj ��oՌ�_��������������'�,�ɉR[8a��F�e��E\Y����b+{�����$�0ٜ����lg�����TLz��U ��U�Q*!ˆt2��K�(��i�(�68X����g`$W�祙m
&���g�}�|�X���=���uD�@�i�t�M�N[�^:�-eq��ۓGD�E� �~�J&��%���
���Y]�������.D�3����{�ǎ�ą����1Eӷ���=4>�ƥ	����s����6���z
E���n�(�̏�I[ ���q��3g����@��~�S.�1H�^�s_Ɣ��=Mq���WI(�� p��$Exa[O`�ң �WD�ӽR�:�D�XR��@�~���p�E�H��	�Nu��m`�ݶ#U=����R���Ʀ�aj)G�3�����SZ��:Xc{'>�r(Fi!�~x�m'��1l�z�X�v'�X\ݒ�F/��B��[+}���^v�����Ӱ�f���U|����,�Hg� �E?��<h����N���ZbB'ԯZ�9��y�K�����~l���0�HQ��]w�<�깕C�Ҷ���2�(���r�+* J��[9�&A��Q�4�'�r���ԣ��D)1 �:�9�h���nȿ�o��=��5djr��7nc����]2��͖Wc����� ��.>��H(�Ü�0	�%�W�>IC��W�`6�������� B�q�G�k���+9��Ĺ�[�D!�����?S#0h���0��hGA�(��%���*��q�x���9�;#���}�q�]�����k��Ɇf��H�x�+*��EߙSÐ�O�r�In���Y������ ��6��M��k�}4�b��,��b��	nU���k�֞!~oh�k.�x�Fi���F9?n�g�^��]t��2J=hc���\���,!hϬ�F�S����(��Ɠ<��Y��+*��&��������~8�zO�E˷^�bX>k��$�e��R���@�<���*|] '�C�ț	A�s��s}]e��R��Rg��p�v6P!&�D\ Ny���'P06E�i��be��|���l��_dM�Ȧ)iW�k	@MߙzU�f*J���0�����>���� �\4���pr��i�Ԉ{ʯ��ӯ�Jd��4�_72�l���g���4�Eg���܆�vЏJ�'{�+�z�C\�x������>�"�:�G^i3�n'ߣ}�>��8�"j����aBt����L[����xHc��5�M�B��kJ��ŧ�*��v��hA��k�4[�r�ݫh�yo�j���h\Tɪ�u�>� �����$�O0]5�;�������A���`>߄ek-�x[��m�;���w���%
�Ð*|ī�x�� ����l�\����<�o�Zk3��%9s�i��c*��F������9���U��2�_C�ǝ��7�����K\u��8l�**��O��x^��� Q)L] �vԿ�$-�I��Y����4"�A��p�G0�3�v�u3h�ê����O�W��Ӭ�O@ᐤ��ثox_6��� ]}>l'|'�{(�7Z@�+�b\�X����|��;�՝k�8�(�ɿOP�i$hN
�H*\�����!��4u�dYl�RcBV���pʇ| ����(�óŬ1�V�.�bag�Sw�,�Y� y��y@�2 W�a���Z|������I���ޣ[k��B�G�X�(���K3^���+p�Q9�A�'C�d��*C2(L~�� 3d�Gy>�x Q�t(4R)�B��Z>@%bQ ��ɞ���
���������{[sLb]�[$K+r��jy-,ړ@���"T.&�x�0�C+����D���*S-���}�=�5i�R<���E�<�����T��ݶ<�2��Lp�a���#��R"�Q�E�+�Ln:{oDn�ɾGT.]��g�!FF�Ϟw�7��Ҳd��^s�����x
H�j\�K�[��=͛��Sd�$�g����E������S�-z[_�|�s���*�FȐ��G��⍮3�$��58�q�>]��vZ�B�jA�PQ��МZ��:k�`�T4W��Z�k����<��(3z07~'�C�I�%�#p������!��<
����A9 ���5�~ � �I���6=_rf}� ��Ϻ{.�G����Q+QW �k瘮k�{���\�/#�j�/�Q͇U�KS�a��>���c�)��S��,�^\Q��",E?�E9w���I�p3�l��擡(�����P�*R����.�j�w��(d:�)�n	L �.8�zz0��l.��qh�Ŋ0鵨����V9�|��,?����gz���.��h� �.��5i�@�?��j�
�8}�gM�<=��Uwz)��?M��TqY{��߬ʹ5���I3�d��T�WAhXI�F�2��P�����dj�{�(���C�ML2���cbj2?cQ��J푳e�e��#�⑋5���DH~�2)c�zP��8.�
=��y|�Z�l�6�ڇ6H\`��2��~d��r�z�ѕ�i�@�/M�����+w���e�!�oz+�k��}���Y�C;��s�bl��M��5�_����6kd��Jb*��4uR����T�U�,h�8� ��V��ɞA�Pފ�T�5�975�Z&^���ڙڗ�)�LIZP|8'���1�}�=���4�ل���;?��w��I�l����}����xQ֔X�[:e����gb����+e�	xX�[�:��Ϫ`.�G��Wj�'w#���v�A���������d{L9+o�&8�ۗ�IB3���9���I��Xj^��)a����;�$X[Y�1?%Zj/Ӡ��S�b�*m��Z���5<G�k����b�r+<�Bh,�~�-Ĩ�Q���֯p<���g熮����P������ю"���yܵ�[�.�i{����/j#�7�:��*yJ������_��xY�[�y2��������� G	����� 6��@�}aql���w�{��dE+(_�Z�J)t���Ν��N"��?]��F��W?b@��RU:�#��:@��_/������, ���T�J&��~�Q�빔����	�A+x7k<���ɛ<^巆f��kq��?�KB�����:pKΎ�i�1����{EJ�L<*�+�.�.p��*r�B/Z���q��kz$@�U��縅(���6��7#�O��.Ǩ�N����C_ɩ��Iy���/bG����g�	��`�U�>�tZɷPD���]�vrw9i<�W d|\��r�Z�^M� �Q|�l���_�`uV\�����ђ��Hi�y��g�<30��sd�?jet}���=��f�/��{q�^��*����]�}7i#�:@=�?�ͮ�˘�(Q�<��D�/�k�����Đ�`���7��<}�������N~L����,�4��"�-�;/�Z��e��#f�+l�YC�ո?�єl���_�~�p0����q9g̝�M�~đW���i,p���*�P�׿[v6w>c�I�o��\���$�cA;���
�3޾�.g����D��g!�)�ݹoԬۀ,G/�Z�K#kB������u�� �Y-�a�c3�R�hI�|�@����x��_�� �,����苹&�m�MھqE��VAڼ�I7,�F��M;?7��'�W::��j9VL?%I~����s���̯d�:ڿ��^��:���-���ʂ��/(=�˔i���\h��
�8Nfr�L�y���f3pB ����_㥰�f�m��2�H��fpl4C�-�_��i%q��U\1G<�>w�b�a[]���RM�=��O���W+TѶ��֬Z�C���U{o~cwҘ�4,J?2�)x*k	T��/_�8��؀���u�P�ʅUY��H�"<�j�Qt�Q�J�������JBپ�X��!W��\-����-?��'7�
O.��>�j4�kXe�8�|���Gc�l�I�H�	+�=��@f�m �*��#��H� ���������دωƟέ�{�#�o�X���L����S�lԣ�}���=�E6����*nz*6�AwO�=66��ھ}��j�ƇODR^}X����w{iim��-%c-O'Ί�.Y_�LH[���.���~̿EY	��S��%�����cqKԴa����m*����jc.���*�lCx�0�	��7Y����Uu��L��a�Aw�o�.]�wC�V�j�CT�#7h}� �o��=�-���v$���k�y�>���u�,�䀲��E���.@)X·}�(�톴���\�҉r��w\蛋�%{�E�BՃ\۲L��1L�J�J~8v�_�3�hچ`ti��KH&�G!Nmv�&J8���#�4��C�&ĊuX�$�A����}���?��	 .4�$��&�J��6 �-Uބ'p}T��T	ʗBl�0��Q6U��95�`F5\�9*���	��(��vQq\���a�T�?��N�MLf�h��Ύ�����ܵ�R�l�:��y$F}����`1@��j���F����T���Ξo�3����ڝ��
����\8��wH������:�[$��krg��
�D�ۍ��E��U�����s��A�@v��@ 8�G����EAa���cG�4-�l�7n��zD��6�s��{P�eI'Պ,�tcd(����Z{��V���?��1��]�f9\" oَ�5QYMrI�}�^d�ƀ-�
����dtXR�?�%�-�%�JZ�HJ<3�`�i�Q� 3�:.e�5���F��,�]cGt�f+`q`�IE <���a%`�_ �O�vsq�IF�O���Aa�bT�Y��_#��Y^^�m��a�z�vϱ�X���(��Sw9s� �7�8���U=�E��� ��z���d:�ۚ������hA���R�)�u����S�S';Nl�pm������m�oX�T����e����!*�v���Qx�fy��L��8��l�pH��q��@��s�\��a��ײȣϧ�0�?Ґ\�t�yܢ>����k�͝�]Fz'���f�K�A�����]_����mnD�wN7�UAy���!Q'G�֏�����O�'y����i�Ja=��.��kH*���j���ά�}����J��F��ۥ)�"?_I�I/�+�/�T;�zaZ�{m:��߬����_����)#���~����a��;ۢ�i/�cI�Gm��[���kO�4��$V��	n�8��S'w�(���}��A�q2ݐ{�/�}�Tra>y���_��t��9�X�g^2"_6��+q�-��fXȢe�>�l H�߆r9QB.8�zl�R��Vp� yr?�R�7���k�Y�l��n���[M�wQ]Be0j2�����'Iv�sA*d��\Hä#+t��u��J:
��1.j����7L�x!�c1�'b�w���?t�����^r���HB2�'��@��ix�R�p�\�މ�Ll�us����!�}9�y�Z�����nt�3U�.����1���L�_놢��\�#l��W�ˊ��敕hf[cui����,s
ƫN ��3�%�Ә%��Mb7�Α�G�	XzzCt�M�Z�roc&�{��Yմ|�*^��t��2��bRm<q"F�(�;q�Rh���B�4}��uc}^���6!%2 9s��? �
� *1&��'I����k�r=���>���'�K�+R_��ڨ��+����ݼ�Tۇ_�k���P��)a�F��|������[rg����v��eV�P�`upQ�"�?����0L�ee�Rpq��vlO���C���2�W2�]P֔>YL9��|���u���NG�<�> �oC��x�H5V�>/FQ�lv���_�n�Jt�}bV5���7q��%4�+�k��y�o,DmX�g���W)U�[ʔ�"-ND2y��뮫���4�k�5��]�v�}z��=���XJ��G���I���yg�_�-
ҭ����YӁ˲F�^b;m�]nr��o�4��'��>J]�	j�ϡ�����e�>�ƨ�~`u:1?�2`)�AR�J����f�ik+�
$��^(�;S ��<ť��Z��M�S*�b�5�.��e�����[ͅi��o�(�H���Ad
O���ZtK{�la�@ښ2��K�H��YS���鼿�R/�_�����s\��߾���q��dV_�]�	X�������6���۬E����KTnX�s�α�*�����%ѐ��(�k5=�c�$n�����
|
ER,�K�@�;F��'�Yvc��ɟ��8R��L~ͩÍ�ӹ�U�M�@;[����Dv�iO2��s�tΆu8F�/�W>�	��c��d�5��'͞�`�h���
b��s=N�k���1?���Y�������(.��!�J"��}`P�H~���L�gj��H���g��_SPS�����a��Z(�����������-�|8�#e��DD��K�*�8I
Mf_� p��X�汖�Nl�iM�����6#�v8�B����m��ʝHDh/L��}�Yd�*��^�B�ɹ얪X�xc6dt�D)���5��,M����˝P��np
���y.�DԷJ-
��_Ԧ(��� ���lJ���{J'�7;	e4�ܮk��5?����/����a��AuT&�p��D��\��	J  �YU����q���l�-�4��(k��]��fb:�i��<(�X]@�H�b^u��o�#�-In����I߀��엎��/��?0��f%����Y�nFQ�Қ,^OX���.f���^+]��n�.m�|"]a�XoR3���X[��X]���G~<n=t9�� �#G��$�s��a�i+}D�?�fۨHn��h���ZO_��L~tg2���=��c��&N5�aR�͛"�*BW�~��	Z�A���!�h'E}#�!�|�i�/9���O��+�(<
��4^��(7�]�0�	0t�X�,AhI\�>�ť<�K(%ÃRA$�Ve�10U����Y�Rsކ�g�s��\�py�ĥ�t}��-���D�2G0Hh ��^��\$t�#ʜ����}�6t35�E�0�� �0�m��Qg���9�s5=��ku��Hh�o8��q_�iҢ( ��5�.����`��4I�!NF=�L'>���9e8���&3�X�#S�ש��m�'gZ�貽̤pb���*H!A��,��}�B���z��芉��t��.,]��D�f��� lyq@��N�Rv?���މ�������yԨfoH�'#�~��x����8Q��#��=x�������%�I�����h�3��SNnH
a�aa�<@&x� -tH=2����dH�Ď�����v7�^�����z�!B� �����"I�>��¯^�����vU�"Q�+�"=r��/�E3��ZǴP~[8H��w�K4�B�Ֆ�/&͂DG�#�>W[
$����x[O�QB�(�ߓ���$*u����9L��z���62$�Asm���]"��(��#����-��m�̾�=\�0�o,
��R5H$
1���\�Sҡ3@-=e�3��ɤ7��'�G "ق���̡q��&u���7OR�U�?��U�t���ǟ����(v' k�6z���df��"U��-6��n�3g��y��"��B\�VV�u�1n9�w{���!~��}y�����a=u߶WQ@�6׺�Mu]����=�2� �p2��t���mh�c�	�'���<���)���ȼ+�ϙ`�-��?\����0t<���¸~L
�uo���g�>t� ���`��< H�̮%�n�?µ���W:6jV��v��	6�I���^^�H��	�03�K)Y�TdxQrDb�L�<��0�|;�-��TR
`�BU^�t)�Oy��?�!���Gmh@�3I�K?�m�o� ��VP f��iO��9�ӥ�w4T��٘�M�+w�	�͒�K$A�4	��8��X�<@�/p(��-�/���`�Z�����Pڌ�>9UUۙ`#|D��z�3L�Z��K�\?�ˌ$�Y�J$��)!etሶ�d��"zy��z#�A��9^��'|�2
�l���������gmas����C<x�\��7-l��*�3�H7�R@]L%�O��6[�R�.ԕ�2��a�w��Z	��'�� ����gH��cтp❊Bcj�����X�����z��r�3�����t^��gW^����A9S��"L�?'��u��<|L}��<�;��L��EF�1ڍul� 2j�S>�3��q�v�1�J��ËM^�?�Q�h�`)o>gƗ���}�c�e��r=ԗ�����x�Xد�^�w�MWv#���B�g}f��� a�2ۿ�ch�A\#��|@��c��R����	�U��|��t�����:;�Xm�#���aRC�b�8]`{��GS�U�_�g��7�0�R�mT袬�Z&�/֏�crGȅ3A�2�i�y�E5-��l�v��N��?e�\�8��M��v|�Ux�a� ��OcBu-�ހ���҃A�m�;��� �P��=  �J�X�2�/U�C�/��6�h8sļ��U��U¯[ �B�W��n���řo�y�'�#T-IFg^�rD�{����9�l��po�~��5#{~����&��Q�	oA �B����2>ա4^m��p������.��dv�uu�'U�W�/$�n��_֓�~ȹN��ԛ&NR@�D?���}C/��ёb�.9gQͼ(��ͥ1�n�������Y��7b��U�]?�XQ��nC79�t�����y���������@l|���A~v1"�?��vݧ�`�^@�V"���7Ѽ��~XT�:-��u�?�C?c̭ڐww����׍"&���5�6��I�����3�$�|���S��'?8�%�z�x~λ�T["�:%^�J��\k��^��!|V�<�Q�*w%�XF?�A��_�'~s����i|�(�8>"6��?s�҅ͦ[7��ЮOr����3�Pd��p%}�L@yB=�4�rs$Ӎ �@i����+��%[�|�����3�~[���k,+%��2��v�Np�ɰq?\�$	�HJ���rK�Q	��	��R�E��~B�A�A�	(:]C��_]�Z�}��2k8GĂ���u�c�Ef
/��� 4��~��P���FEs��r�k'v��EG��O���5�I��F�駛�ĳ�a��P�SC�׻
�'�g���HӁ)_�iq�s��>�$E�S.�X
��  �;	�ZI�� ��F��v �T��Q��ɭrn|�7��7�
�V�Љ�w9=�se�:nPr�f���B�ʾe�/�x<�A�	���逕W^K�{��>��m��#�豳�-������M:Tv*F�k��n��Q��.hc<as��$+����u��,(+����*��T��o���W �Ǖ�l�=ܔ�VM�����7������r���Q]*e�8-���̯�	\��Ĥ�q�%�$�������"�jQ@^a�|Cg�߲�w���&�Hv��fA/� �a�S��г27�܎�:���<j�-,m��*��*4��!Ĳ��$���%��j̼�.,���(9��b7�/��yRh�	�P<>��<D%���9z�},��#yػt�Ŀ7�&Y�[q�*D���@c�/_ˆ��~�P 	8�n�%#�		����WS��a�Ԡ��/�Хp��"{;�[?v���dg���ܰ�nl�]�x*���/����!��J�{P��]�JGX
2��nb�����D��(��XQ1��R|c0]4=�8WVU��n��g%R1a�g�Xd�T����&��@셏k��e�쭥�L����)��O]!B�u	���/�ˀ���������d�x�LƋ@�`ۇs?�u�[�^�$��T�T>X����dr*k�ۛU�tO�/ ���䷙V� �HK��<�_�٩־�EBCn)&/��m�ػ��('ޣ2�v�N��^�4�Nj4�\�;\#��G��a�N� ��d;���1}(*��ٹk#	f�"�X$��^���-�dI�u���80�`��aV4֐EL�F����G��5Ϗ~ds҆�*��AA$�V��2O\\M�d�M���7e%#�4�@4�X�ERQ�������_Ps,ōCt$�M����*g;�{0�f=� �[��91
�^���
�-�.%�'U�P�yr����;�C"��k��$x�5�xw�����b]���s��9���E��MnD?��B~h�_%ĆA`~-mW��W���E�0~#�F��~��}B1����'�¬k>�S4�T����Ft��ke9��G=#+� ����X�gա�<���t#\	�O�w�]�����ܘV�s7`U6+2�aǅ������v8Q��
��*�;�0֬^	/Ԗ�P����;E��+r�4�L���=#��N���q%q�b�O�ݘ��>�%Y�<�Qa���2�xP����g���fy�V�}��-�@`G,p���]�3��u p��b<�/v�]-~=�i=fR��m����?�y|j�x�W�Dʫ��Ox��"d��۵��H��E�������g�=�{K��i/���������Ȭ~�#P��m�w��o�~T���K
���>�� qFS�@|zE��	1��W�8)�>��(����m�$kK�����c���6N��9���q\Θ��t:�9ѷ�_8��T���b2 �h+A��w�bb�%H�}su�O�i���UK���s�l��H��lƋ��h/r�O����Jr��Zc܌+���|fD�D�%`F���i�c�Ѭ�Se�,@�o(��d��I+sfJ0X.���Sȫ����HY	%�h�08H�5V3X�#��ou{��cʥ=>�'���.&�k͂&��f�4�f�nu���um��ѭ�����oh(X�n�K^��.Ԥ��B�
'yjj;(�[u�qPɝ,<|��j�	f_��&7�Fʸf�����C�EP�7a��Y���LJ��� -�\]a�?\�%i�.��ݛ`v���(�tq�;B�"^M ����bt8R�3OiVQg����߫3bL
��>���2�g~�����A=l+-Q� (��aeǻ?�mƔi�Ģ�%h�w0zYGr-2m4���vJ�삉����W³��	�6�3d(�@;\m..u9�d�A�Z�5D�^H���U
,�p��o��*y�M{���s��
�+�	à���Gq���ň
�O�����s�Lb���j�8M�0r��a����2��՝��8Ǣ�\M�#~XxC�#>�GI��Ӫ��m��w"Ȧ�WQ<�|"Lz���s�6�����G�pܫnN�͎���سR<�L1�bKmĄ�V7J�f8Q%�Ku7S�N_�L*��2�/l*Oc(�pf��Ա�!�|�i�+N�@�?͖�i �,'G��K9u$���2�"Zv�"�2,�n�����u&p�R?�\m�S�%#0I�J������^���|�>���A�ҜTa)���A�� ���¿��yLݤ_ �Y8���AJ�Y��'qg?�|��a�uA�2G���5�]�s�t3��m�ǊZ�w��;k���Q��(D~��hփ'�\�❻L�_-��k2S����� �#tIՔ�`��p]�B[d�*-J�DUEM�+���m@�0E{�7ԝ�o��V�Nv{�O�wVxdX�@�b܁*�� �+ax�A)(�]�gY���!��߅"l�h�[��K�j�p߳��vk �*�y�ƭ�ndY���Z�U?'8>+��T��Ɍ�M�*����h����s���a�Y��'�g�U.�908����՟[[;���}�FQ#�蕐5rߏ�=L��|7"�#�Ѹ�6���U���-IT��]��&�LW�̀���~|pd�;�cQ�r�nڴ�5K�򠧌�����YEEvmH[���D�GW�:�h���y�A[���R,5L�����Jb��
���󣶠�Bp���<@T\T�G�Ϯ�j�%V�Y6|n!�,$���ɋ"��gd�ёRg���dh�;21�|�Am'Iư�$D�@s���B{Ȧ�;�e��\k�����T�'!��Ü?w�ƉmC����?�k2�����Nun�NkV��n�w�Q3_����S��Co]ԫMuHi�iЦ�Ć�$���S]�B�n��ȋX��&�7�/�?md1�Q�"E
�U��:�5�bx$9�6�<'�E�	"����RF$M�D]�t���Rʑ>�9<��	�T�����5Y�5��F;��7M��e��I�P���W�3\/UW7�Ɋ���얋'G�(�w����%z=��+�>#%�[���n<�1�{_�mP��S��B�*��Vt�.�a������7��I7�$�L�bjc"�t�ڠBMz%����o��eZ���7��}S��<���/b!�Z�����k:)�*��h�[���2��J��f��Qsz%�F�1I��@Ţ��9w���LCI�I�Ɏ��f�҅Z1����_�#U?S	T�۹'-O��B���f]8����� ��'�k܈Boݧ���ݒB���Q:$RW%�������q��jM�s��(vŐp��0[���8��RWN .?Y�7s�Uv)�Q��~����R�]ʉT�>������I��~UYG:iMg~�W��i�j��=Ǟw�}t��������x�J�Xo��[�tS(����Z��ݓtD��	>�c*	rH̍���^ÄE%j�Gx��(i:�{*�s�+\�&ƕ�,�d�͞^��>.��qǓ�N =EΏd['}�+	"�C�!�T�k�RML��*%{a�%@��$��`0
�0d�����uK��Qܟ����W�����4L5��җ�U�V�)X�Vk�X��\c�l(���
�@�@��I����)n�mz'���B�A�@^��Bc���h��N���h}A۟��ɛ-�I�C�m���ʫ����������|/��"O)���x�m�� /\*��E���j����=H�wc�O�c�:�H��š��]ǤOg')'7x��|"�Q<���G0�*�.��`��R����ĕ�l�l���a:h�)���2v�fp���}A-K�@I�L�:�d�ۿwůi���m�@,����j���=����_�?�~�q��8B~�H��L�ɒ���bb.s��,�o�u^W5ֆ��T�����,�t�V,��,!#���g`��Pn�1��ݦn���,���̋۾�xv����g~2/���ə�5TԬ:�+���9[���.P���5:ިP��o|���m�)&�H$���j�'�3�S��lh,����0�>��2UeeBG>7������Ϭ�́�Zk"�����D*G�z;DЗ�0�I.��ŋM��uh"m�^@	A�Pͦ��X�ːk)��������Q� '����<{�(��qB)O�<�����Hȱ��Rw�t����PƖ�p�?���@��"�zs���{�!���ŷqC����hh��T�)�]��������9��O�-��U}��kx�.,�*[:�v�$���7��dx�jc��"����3��<��Q�.�>6�᪟2@$��?h�9O��M�q�&�@�\i֢��?��������s�s�q�
@T�q���ϵ�ai6�?�آ-�����Rik����ܕ�5����ƝmZ*�-��q�����hU?%k��7��/��t��XD��5����d��Oy�i�Or �k�� R���tQ�����2w�@#���dR�8p�ѯ�\s�� Ë�m>�&V��\���H� @@�B����l�?Ǡ���Rv�5�L,Z��e�#�',n
l�W���EV��B�Z'T;��G�/��$���m������	@��PH�Fi 7���H��y����Q4�)��l���rZS�iX���5'�h�s?KY��W.n�a��O,!6���9�9�r�	���,z6�n>vC�׃��ꢳ��N�)I��ec:�W�X��4�)�<CI�fIyo�vn�у?��}d�+�r��<X��a�%��T�P�"!;bٔ���j�#�Ϙ������lڴPޯ�Ao�|�1���uE=�R:#_
ɯ3j�5g���������2�Φ8
��L7]}�NC���u�gaN�����?���Le�$�ur������:)	'�_r[:Oq����@�� ��v��5�V�I/!K����7	�v97k�b��V��g�/ܪt]�* �a� ���x�5�\7���A4&4�wέ���h��񸏿��N?�3v06�~�����?1��s�m�  �1s��<���7Ր ��p�A?��Щ/Fʻ����Mبq	�@�%����	��R�� ��\Q�
	C�'T�<a`�45"6J�G�?J�1�=��O�R�-�qe��j�W{�x��T
7(��<޼�U9�R26���n���ݴ)�z+��*�(��w���%��$��98i�O�Y6�D5��[��IE-��b�V�`��bH�:˭�f�JdV����.Lx�;@��j�qj2�|^�:n��X,�#���^��V*؛�p��NV���� �+SG"I��E�z���$��aX��m����:���=�3�q�C[�l�lup��@L�o�7e�8 n��{�.�o�Sej�D��j���+��u�azoi����%w4d8LZ�	�S�s��p�q����}��G�S"6
�~�u����M�$N�q�M[�c��o	��v��'�G곸V�~�@�iғ���p=&�U��m�&�S�[��v8�_����yf��gT��?�Q�m�$&`��;g7���$��p:�=�D�ݍ"�+J)����H��1}�I�g	
�O��ŪwƊ�{�t\�{�N��iC�FX�@��r�t U|ǈ��[t��~.l�^\
^�&�Z���؊���)���7~���@�]�|H�r�5���2��lf;B1�tbG��sA�\�DQK��3�q�_P��_�v5-v�$2�HUX�o�t
�(ad.&R��R"����7���>TVu�\�J����7^8>q|ө?��tba�����K�ލ��G���t��R?L����R��6�f;�=Ζ*�� f�P���P��
��1>����6zBKyE�{���}y��'z�(�[,���.͹y�Lˍ�����X�4����WW���`��'eQn&�>>̋�'/~�n�A^��0�7߲�G4��r��,�� ��Nl��|,��\�)��H5���G�f�͊��X�U�TCV�6XE7�O53��FhG����Qb>��� �����ә0�1��p~\+��U�<Eִ/"{��kDB��*}nR	��&�'���G�s��o��?�	���"��/��M�x��nwE��##�G��5X+l3��j/X�M�)7Uϓ�w>���B����i2bv6}�����fūF�E���gˢ��k���L��
((�Tso�	�#�?��F�<�rNz�¸�6Wp'�L&J����Z5�0�n���Q��C��je.�A�*����~��� D`Q�K�:���7�呋�����OOH6�-������f��8d��C��&��GA0MmD��mkK�4ı�utPbV��$XiH j���Ԗ4ט��ٟ�Ȑ(��=Y�Gp+_Γt�ܑ>Z���V,w���K��,��»0]�ͧ��Ѱ����:b��q[� 0�y���
l�mYE�p���|`
='G%#�!誤�-.)�O�A�s��ďG�k�9�*QҤ$��"+��2�b`��W8rե�l��9j�u���l���.c,A �c�)k
o_>$^�4LyF�k?�L�l������(���`�^��7���Z�bWt�,!���;�Q\c�O�"n��j|�<�9*�����S�{�V&��SuI8�����x��2�i�X
C��ǾA�a *x	-h;�4e1Q+��JVvÀӒ�_WI��H)�m9a�~"siHA����N{�K؀z�7�jI,|��i������2.{l�n����W,?�)n��o �J��=��Z��b?;���ݏ�WQ٣�QAv��f6E�±���N
8��e�H6X ����e"�Z��=�h%�>T[�Ɩ�zF��=L�&�Q�|g2[VK��nP0ҷC