
module debug1 (
	probe);	

	input	[3:0]	probe;
endmodule
