
module DEBUG (
	probe);	

	input	[0:0]	probe;
endmodule
