��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;������D�ۿ{'�����`���T!~B�YO#G�hE��xqd�l��O�����vi���C�x��y�Zn�Z
?� ��w���`1FQyb
���&�8�Q��]�
q?�O��;���%���Jٿ2ť�E8���Xͷj�;�v������Q������9��Y����s�����B��&��+&�L�\_�9Ʒ��"�H��1�_W��F�����P��:����?�%���=�0dù�e�Ic�\�􅤥1Nʟ����U2�?7 ��L�Y�{��5w��gx��o��E"����
��+�!u��g�6�2�,n*Fv��AS���	%��cu����b��M,�
/�U9��~�SaT9�m�'	HFǿ����Ej�o��L�W~ � ���ɑ��=.��S��� \ �of h$J^\�u���qQ�'
A�'�w�xޕ`���ՇD�G8�|YD���=���jʚ�s�򋀠\ӡ��o|�:V�v�\�c1�_�ֈ��s��
q�"sKR��Vn�مa�zgZ/�KP�¯�e&���թ���\�p��4|HKw���90e/.��j�U���~�&�H���v�c�/!���x���D��JM� �C�� ᖆ�l�X�{�sd�
�w����΋��E��~V+�n��R9��k�έW{��=���q�?�a�m��:?��V���\�G����^M�"�{}j���p�7R+���pEȷ�BWN��f�J��X+��S[r�����(�d�+0� Og��B���Ϫ�-.��#��mm��}aV�X������&[� e���|�9�b$^�&�j��Ķ��oL�)��X.(.��Uڡ��!�uH�a!�RP���k����?'�"�ɗ4�;n��t�k�@c�������f���'�,������D`��7�,��j�WOF�)U���o�/�����I���#V�G��P��[��l�e�GL�"��4D�E��^+��3E(sh���E��x��K�H�lG.'弃z.{#i��o�4b=�]�����S��M��1SeX�� ə�ʘU ���@D'��K�� �T��B�=��>��x!4�9?S����S>+�&��F�N���I��P��%��-��UDu� �?|�V����.���K�vԵi�5��@$��MB���m-gb�B^�)���S�z"w����3�h\{��R�tV)�:�p=-������!��
��OJ��6����pOEz�ޟ��5N���2����`�;��]:�_!6�J��~C>I)�ץP{���yڤ�f�������i�Jnj�4�N�'H�(�I'Kie��X�E"���0����ϙ�S�\e҄��_!_*��
��&�/fd=���19
��ds�����(���OS�Y+n�p�&d��Z&�Mu�ySc�>c��eP$�g�a�)m����N��? Kb����7?C����_& ���%���$�8���։�15���/[ڮG�q�-��*/=0L��{kR��S�#���)|�L�� �6���c�P�\�����?�e*.CL��=R��MO�Cx����Q_�~Ȟ�>�.��K�X���q��vv�L_�uI|�:��e��4zD���+m�.¥T�r�E�� �e��#�F���#U^D!��������e��s�hkf͋9Y��;f�p����g6��t~VkɽډX�[ܼa �aɢt4��vX�}����ߒg�=�����3gD�P�}H Q�%�y
	�Q��U�IV��h�#��k.[B�A�����j�k�n-���JL�]q�$u�N�>���N�?�\'7�ؠ}���UA�;Jp
�<���0.L���w=S][�o���cH���T��@�̟[0��I��x�'�Z��o�	 A%�_��Z�3��<��
�b�E��rc�m��>����c�IҨ�^n(7��+�}9�'RG���8���J2_�VQ�;��5�+4ؒ�i>!SD+�b�R1)<���D�C��7|���"|���$�s�[�@��.����f!X��[Ś1���0	J�h]pS�R�Q�l�����j�w̖I� m�l��e 	�9��X\��y��U*#�a� ���.2�_���k�]P�hj���+���i��)����<���<[�7�9Dʳ�Ώ!���4հx����t2�L�Pk"��!{�bQ\R�3]Y'ZV��T��H±4���,S��^]�3Cv�JJa8%q5�օ'p�k��)��/P+c�����;nQ����n�����;�Q������A�j"v"M���,Gcm�s����b��<z�w��PF9E�ҟ=Rqv�m�
Ұu��k�q?�-赘�@���鶵@��~%��މ߮����]�f�ܓ]<�-�$�eM��6u���c@m�?���q�W퐄F������L�+��0d�%1���j2<_!�������=�<��}8DN�̽�XU	��n�����B�\oƚ��+9M'CL���ﭺ!�S�!�k��U>KP�)9�(ė��A��x݊�����Ws���ƚZӧegZo$���T(���v�t4�����a�?jl�#�������:�@���9w�w��g� ��3�U�7�o����V0-����_?@�BG�˰q�xk�$��*�M%�g�1��8�إe���X��d_��&�]���\P�@��%!h�L�ò��C".�L�@�|���ھ��MU%���.�jW�� ��|2$�K�q�%�㣽	Z�.�&����hzcw����# �,����ߕ�,�?!� ��_¦ƍGZ��6Π3L��� ���6a\��8�?� �_�OlvjCu�}���0`j�p��эps��@�*���Di+����-��<���5u���y�JU��hp�8)�Ѻ�ŧa�+O�`�����O�6DC8�9�Z������3YO�<HB��N��s,���
�����V��ߢ�U��4�yq���r�H�E���2��Е�g����r���H蹾��TniM�P�� �j[���Q�A�ͬ��iJ1�9��� �.PN �#a��BF~:Ef���u�Jf +ț���y�]���y��N/�9�&��&�ӿ��/�f�+�����*�溅!d}(㔎:���(���4��F��,RO/la���7]⍕���@�2�wGs�%fR0ph�f�"�1��&G��[.�b���=�&�	~{j߸	#�d	�jɑF�� �\��A������R��b�V����b�C������_�-f��ς�����/sE�{����Ҁ�%�5�"�i��"����6D�1����6|�]F�����n�H5��<�t��(���J��Q�	��,=�8n#P27�0Ҝ�u��$r���i=G�i�O{棡�H�u���w����N��@9��l���ļ+h+P���r+/~A�bS��'Ep��f��#l��z7�����C^���:l͜!�B7�×����}�����s��� �i��Uo
���a`�-�QC�i.�s�䐩�T(�Y�Fۃ��YEo�lp�I�	�/��r�k���$-_q��ɟJ�F�>���8�(}�
�/7u�f�*N�Kb6�S	$�2n�C�iF�%gJt2?�<'tu)"�����a��Q?�`:<��_(IKѯs�wm(/���%}.$_$���$��g��Zs;y���
��,��}BZՎڱp��U�����]M�|��36�9j�j�Ms!��ă|�����($�i+���WD��6h*���Q@�}Z�?�Z�ꌎ`*���+�^���K��1r�(t�A��:z�Y��u�����cTDE�IfU}W[��r&�~�	wW��-�����g���w���;����3��'�q���g;3�}���Q�(�j[�S���c�!�����?�)=N�)�\�(� �]��9�kWj-�gu��Yo�|T��ڡ$$%���iJ� #:��w��ʝL�ԅ��܎'J�l���`����AE��41�#R�P��tX-���x��(u;H�~�ي"��ַ�C1��4rtqz��G�iL|��F�SK�I���]i<^�P���HV����2�V]FF�Im���0���W��^Sg�k� �M��m�p�Z��e�L�6���ȢF���c�%���Ƥ9?�����\Rxt'��^�E�GP�R �aVYg�i��nQ:��]���o��`.?�L�i�2<�%q���!
3r/F�Sb��]�}��c�D$��iS�r����Fu�����Q�!G
�%��P!�����_6˭�`ڢ��l��h{�i*��7���P���r��/�Q�?�EZ�TL�.;<��>�a�y�U�팩�/B )�"%'�Pr�|T�%�~cH���`�f'NUc]�ng7JT/�#xW��D��@)�e����'�NvE�{-�(�6~=�T�6󾷛O�����R����A�Ӂ���*D޵�xy��\�;J�h��8D��ɿǴQ�(vj�˽b�TxWa�d���Q���eªe�uS�Q�v�¦j^�'��'3N�-Q{r17x����f��'�|�F�����Dm������w�N�HFa"���_"�ĢBr�X�b,I.���A`���]t�.�"Mi���r������n�{aX6�P_@���o�� �]�ٻ������q���T�:�ʃe[)�mcv��5RDi�,�=��Ʊ\3T���W�h�פ�^ 2��M̊�Sxd���U$kݐM�U��\��0��8y.0M��b�ST,�]@�Xn �v`�BS�)�'�nF).:�e���\�se�j6��7t��W�������wt�x^��݃���s�w�P�̭kWbVPE����faT��z�<�?��ST�"�-��m@��ﮜ�j�N\fՓ�V�.�[�+���ݦD(�l���K���{��8�eb�˫'L�>�"�-�N�**�k5�3�#��V/��a��4�K�]��tm�6F45���ɬ^H9�h}��\��Ѽ��Z��Ъ����E��(�)���2�S���m��+aN���,�OPܞ�w�O�e�٣k�bf,ܘ�|�ʧ��E=F�\D�_q��|d/Y {�̆S�.����c7�6��Wu�A��vM[,�L%�h�@/I�EZ�s	�L���8߇���������T<=ɒFXb�ؽw�N½�����4A���P�] ^��*>m���$T�f���T�����)����W�E�����ww}�����2u<���^ho��Ϥq�'>���_l�w���+��:J�.A�Ź�_�d�0�i2��1� m�Q�����ՙ��.�8�E�� '%�\�k�x�Ȥ#��\5F�)�-�z��4�)�:Db�(�P��ɒTA*�h6��p,g䤲W�J��.���*�4:w0������vBL��؟��wT�~�0�c�����������w �Iy�N����k��O[�G�w16�ЎN=�qN�c���$ٱ����Y�B��hW�%�T%2u՛���Dy����6��!��������Lǎs΢��˾��0�}6��ω��1Idu�}�%�v����[uC��y|o	�'����k�" Kh�[&y�o�U��.�c>��H���ݵ����X�Ef9T�xV#+�]�hq���f:�yq��d��h�
�lSf�����F�+U��0��3|�X���=GTr��vh~8¬��Jey�XS��$���)(��S�`A�B�1��'Sc��6d9�yV
~�V��d�����-m�-vN�/�~j�����z�@���u�o��ao��4��3p��,^��?R�U}o��Q� ̑_�8����);!\�e?���v_fP�$ �u���d��I@d�T}�>��xV2�ý�8&�6YkKK�N򦺱���1�w���2�&���������	S�ߑ2$5)b��O{��L�dq/T���^���O�������7*�^8sZz��:��#[����k/ԁ��JH��zUZv�YyF��w��]��i�o{c^���&�����t y1��_&9�X���+�}0*�G(ۙ�4�۸6m�����<����#��a�Z�����	�XhG#�CHLC;-�Ȭ��&�|v-/:�<�<5�WbL�����I�:���Gm�jk#�T�!^EF�A7H%ȵ*v���/?�P��\M"�Շ��x����<_��*MI�J��ܨB_;*?��2ov+��J �o+���&X�l��N�{Ƃ��i����,�7�`ɣ�v�*,×o[s�'cp�2u%���g{�,�;W���DO�W�
)
�-"��i�)�v`oyĒ�z3DF�o�]�WaV*Z�nʔ�荚�9�>Ԝ�*A�]���Ul��c'D.��/��s�V1p��2���[w�:�.�5F��2���Z-��1����ZŅ�[{W��(V�s��P4��������V�7L�RA+��P�gנ��Mluz��%`������@���c��+�D�dS\�̄
�CM�7>6d�<4�Qr���4��I��#j8u�&�͗~߻2~ٞ,����6�t+,���A=�R��#�[��������Tut�|��o7�W#i�iDA���(�������j��r�����H�i��h�2��!H״At�F>bs=m1�5	�p�W�b �3��p��Zӹ�%>PA��R ZHEj
�S+�.�}����g��^Wxk�XG��x��( `�ײG�/�6Y~��|�F%ڭA�1�}JAz�hI���-�~�f8��4�*����XV���h�Ff>1����{��YZ��#�i��3.���YS~P���*��}�SH5{Y��ӌ�S������#	��L�\���� ���yL�% !:\m��O�e������I^χ_��慜K��+5��ew�Jsx���jS�0cI(��br�/�_����B���u�p��֦�C�܅q��i�wm�H�Y�f��/Я,����)�5u��O�����m�J���/$�)��k�@�����΢�%��Q��D;Y���z>��GQ��&��_���V�rר���IV�ӇI^(�;푇���D�8���,Jlq2���}��`�~Z��I�s�<\������uY�PH���|�����Gz4��m���x�+��'�j�T�!LAɿ]�4t�"�fI��Ƭ^�(��	�`���VU<q%Q�A5Z�ȷ��s�kmN���q�m��m�8x��I.��e��ٗv���mc]I�d��;FWփ��W1�y�ߧVPrtE�daw=v���z� �v<$~�z��.}O�"��K,���Utc'���dc�A�Pf�ٍ,��e�����.#z%�^�H_D�ћ�\؞��ڱL�2�����,�{��WIh}$�s���ZQ-��`�LI-Gr�X���߉���g��"	�����,�RⱉҠcv�q�>]C�wt�̹o�Òof��FGg�0C���)�̋���{b`Ph[����0dn�F����yNÂ!^j��o�ґ�� ���W(�	�wp1Тm�3u
$%��S�4s���m�K颃��Y�[%2��@�
@!�[.�p>��J�J꺞u�%M�Ν&����������Eʹ'�粠q�t�1 J���cޤϬAeB�8^&����}6�U=O��;���!�\F�VM����Q��&���zh���$�\@ױr�	�_L��ۄwɶC��W�	��r���F�J�*I�MK�'�Ry���]��3��V���[q�����.iq��q�k5��]�rK2JmO�b�Z��oan����?�n�~a)r�+_hs��Z�����9K%���]l�	�i+�����H�������	������L����~B5�:~���v�����#�􇴇C��u�RL�����[���72��vw��>��"E/&2|����~��z6��&�jW�u������ï��8e������X�S�3��ș���rA��\���+�F�ӏ��?.��ɾs&�,d�c|廹l��ws'��lCR��i�Ze���NX���.?RRZ@st������U�X���Cs<љ)��T�(�f~�8��MX���x�_еh��:',F��r�-�`C���o��ɭN�G�jefH0A+O�#h�#6��/2�F��p$tY���t�G'S̓%�[�E<�3�ЗR�՚V��
�3G�k�����%�-�{����*%7ޕ����������N����P,�I���H�b����F���$��f�	}�<��8eh7j+A�.����昑��WQ���4�@���5m�	���@�B�m����w��x�!�mP���F
,⢽�3geg�I:��9[w�؆���P*ۋ�]5�v�niܟ��n�L�B�����G���gk�܉�Q��Ǟ<b]yAS��{G�x��2�����銖l�#���Qo����a�b1D�9T3C��@Z�t@ß2lېq'�7�1�-��sX���L��/�檝t6�gГ� ^
J�ޏ4� Z���l�j��������+�lC�(��GY���{1y�
g;ɟx_@P`2 ��G�J9�ZZ�$%On]M�����*���ͯK�o�����S)��PwK�0���,��,�;��3ׁ��g������x�e5��'��xS�IK�<�k��(Ȋ��}�����1x�5��*�����O��C]��l*�n Ʒ?���chv��n,�� �cB8B>r�vG�5a�����3������]�e�d�f׌��\ Q`Ĥ�� !:aͥ���/$=��=-�m�Q��/� CW�����ۄuo�:! ��഑��Ϛq��$a�:��96��U���"��x���r��ހ���څT{�6u,���/	Y;7Sn;�����d�z�V����;}��v�{����Cz1o��=��R�La蒕�G�U"�YV�CS��[o��!��D�h��G$�^�nsuf&�@�/!�џ_ռ���N�7����L���'%�y%Me��H,�>uE������\���N+I���lo�ߕ���(~C����RA�>v,�J�F1v�����?�ŕ���*H[Jí�t������j�`uR��66������.��hne��A��|jJ��R���l����҄x�&a3;�߮8�:&�C߸2~���u ��(���Vx����0�R�wA�7�5:�>O����gx.�N����@��-��_��)Mب9�="�n���aF?Y)�T��@�� �S�	������������$iȓ�`j��&'d6��#�d,��;�sn�4�@�=%N&���Jn�q^�v������&� 5�v�?:L�Ҩ�̍�@�!3�j��˱^A_ ~�&��bdo!C��z�Oqy?�q�`*J���ANh�R��gn*�:�> ��Ak\l���g����Ih՟�%�"��A��{+Ӿw(LH�+9��w��FG:�*�DB �(���.�(����ԬH}�HA�Ik��lކ��m��� o�QKS������`����e�F���֙�6���Ikb��[~� �4i�ő��E6az\�B+GS�Lk��M��s%���j�V�?f�с�h�XBz��Q�|��Idt2lg̥2�u��$(ǡ���e��o�H�1F�GOP�b H�B�>�@$k��ա�=Q���^�]�>5���}�]��H��BE��1]~M*xz�J�0�w��N����r��#�f7.�>y�I|�r��:j��w���V�<���^%�	���e�nLc ȟNX�u�{zs�
��*��6&���a.$.df�(�_��ܞ��$����Lޯa��1"7�E@��)�Z��V-�t74$T =E2w�\�4j�h2P��ę�6��x�����c��8�'�ۙ��L���v�tF�?	`��c �wTa�9�j�ת���/Ŵ�!����ȟ#�.;@��K4�v�~�R��/�����NZ�d��!,F](
������ME'u�=*��AȬZ$�S ��f�`��_��U1���s���E&������ez�|�Oo:������Q|�h��8��� �&~b�[O���L=�:�U�#U#���j1���n0oз���9�F�R+� IC���#���#��<�@��Hc񦢱��B�������:��fc4�fӓ��1��e���<�)��N3?ґ�z���)�C�����!Qd�����	�?���J����p$N���U>4<��hxM3�;�O@-���
b�  ),�)\IM]:R�`]����>ꦭ`����r�R�s�����\��Ĺ��_� �N)�sdtA�ȉ��(��n`���ϴ���ħ�ڄ�I4o[{�h�W�61u��!���8��4)�΍�E�=�-LfSj�=Ӿ ��1ٱ3|���JX>Y���TJ3�9'����B؂���2���}��j��E/gh���Q_�O���{cV0�:�b��a�Q�l�`э0�9��t�/����ZA\��"_Y�.Z}D��^��e{٢p��ð_X��h�J[�,l����y
�aO��JK��E*Z�[�3���+�pSg����h!���e���Dh��a�du��o*\r�$�Fn���su�HA��]���a���/�p��)��,�H��7��?��egX#}��4_ʽ������+���vQ�k�}у K,j��4�د;1{�a�v�$�w��O~\OI�`>�V�#*��+�^��N5sqru��*શ���.<�k���Q����F�	���3���l}1�����˱!�o�$�k�JA�N�qe0K{�-��)�����=X�Dg����C2j�^�:��m4�Kl����?j:Y=�K?���ճM�':@2ԅ�*|�%-��v|����)�}|�Za ����Q-�,�{=��������a�3�.yH�>�r1Ʊ�`&+�5��NɾW��'��������)C��uX�48/j�7�&++'[����S�&��tk��VZ[�|����������I�����4�1���
���4HH������\R��f���!OrFYM�M���ĉ�ؼZ�E������mD�����5�~�N��8�Z*��X0ʙV��I�X��c�F]�����r:k{��S�c8�z�g[<�m���PV��a%��T`��e9WBT��K��(��A�����[4-���\�УmYZ�Kq�O,�;�����qW��.ZGeZ0���B�Ɏ4:C2�ąˋ˛ڟp¯j<�]\'k��RU<���F�r9�l��T���A��U��!�D�L32G$���I���_�0�Tn����!���{��|���� ol�5�H# �8>�/�/�,A�b5'����8���x	mP�H2��જ��N����$ײ��Ī:܅�MՐ����h�B��R��FL[	��q�Ɯ�l�����Z�^Zʅ�Z��ã�$5P�v_��]z�#�I��������/��plBXS�
%#*��xQ����)G����=ⶼ�5A2,��GՕ\;c�&��rP�(%�N�����O!�]v$��t�����s��Ov���a�q�+��'qD�v�ϙgɬI�����B�;k�X��"�ѷ�w�V#xH������{�޳#�:�d���Fs?5(�[�<Z�0��_1sA)�m҂tHҿ3_Wn8[��+�2��;CF��]- ��7C4�(�:�������h+\ĔU�+6)����#M� ���"���IN�����Z4�������W�uy��aYU��3w��(�HYߖ�b�93j��
�E)�;8.j��>*���6�������Υ���7�;{:�9S�-~�@U60T�o}$c��n�v�k@'B(�F�XE���
hE`?r�侵-,L<��Dj�R*%�C�Tx��R�����ڠ[9�q���8rPЌ2�`��P)e�싍j�q u����v(�M��3�(j�=,ċZ��N^!��´5Y[�Tq⮼�C)�7��s�O�?�_7i2Z1���H6�%cM#�jz��e��e��o���ۈt[�����t�w��� �\2P�2^��I��w�FQ�?��}���o��PCx�k�E]�3)w��N#�"�B��M0ƾ]U[-��i��5�Xc]ο��e�0��rC����xAژl��ͨ� ���5��(��NԊ[�u'�#��w�X�M~G�w�9������{��60k��v�% 6�f:����sh�ۈ@;�%�^͟�kg�d���I�|w��S�Z*z�.�U#�8���DC�����z�*J_�vT}
�X������vb��x)�ѷ���b��I��2m��c!��[�{?�S+x�,���'��$~=Y]�K�ր��`x%:c��7��g�Mи2��g�����0$���9�T8eq���hJ��=C�)p�ND��B�m��k���z\$hYܔ1��?��'�r'�/��J�ȗ��\��Z��5�J�&�]��