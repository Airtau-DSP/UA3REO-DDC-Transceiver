
module DEBUG (
	probe);	

	input	[13:0]	probe;
endmodule
