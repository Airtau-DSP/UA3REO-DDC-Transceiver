��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����թTgQyQ���4�.�7�,����R��)�]�����博����iad�.Wh�Llx�@xgb�WQ̓E�-A[��6�y������cnD<��0dJ�ѱ�.����p5^���A�*i���=H|Z����ʢ�c9ʘ;n�1���=�(��`�Sn��><.D���E�;3���/�Cj|�(DK-OuB�Џ_�k\��,��[ �����i"��N������nl�c}`&�xS� <�g�8D>�K�M&�횮�g�����i��Ω���a�S�\fDf�?�vBD�fK���5N��;,>
��3xg=e$Ո�1�[�Jà����k����Mel!Tq
��{<z��_��F�����'�w#���J��Y<X }HZ���f�1��u���O��8�k�i��=�趫d���K���+/�哅,-�_�a��Ps�]Wy5uȵ��� ��L+#�����Wϟݕ��b�}�[|_m3�:�O`�ɖU���Fj�Y�$f�f�Ɖ�Z�ľD�S2�ߵ�#�w�i{��������r��*��]���?��/eRR��~��{�l��.�H��wpN�!Sv��4��ܠ�,�"�lE�Ǝ�(���g"	6Y8��qW�'�<�>߮��:q7�݃�D-'y��x��
�� ��Y$��F��g�Ij��-���rv*�6V���5O����n����ˀy_���}��T���Aþ�W��7RM�V�8��!.P�)e��>�Q`,UY��>~K��&:<��#�>C�5�w��)@	���sM��J5�"3� �Ʊ􌎌�WT���5��nږ�	�JХt��&�/ē�o�^"�-�-/ @P(<7�����nG�4���F	�%�Qc�z�� h��ul����ok��\�(J�y��S��S;�S���o�嗍�Pڳ�W�cȓ� �D�V���MD���,����v?�h�FF.����Zǖ�Q��@��m�cY�͵���1N��U�c:K �#NÃ��)/7E�%���W�Kı����:(�L�R�Uҍ6r>�+�z�]-��)��\��X���ʲ�oJ��P9��=>�C�@)��P���VT�I�C�����v�2Ö];fu0E_M�}�n�ąE��t�eIQ�|�a�y }��b�@���̤�=�ȟA���u��}juE?y�b�=�;��ҟn!��ⲝ!	����  �&���wdz�C�Tg���ub��>T��(B�B�Iy��<���o��]}2�@��@��PnC�v[,�T������(ϰ_����G������"E�D�3�+�`f��םR�5f�թ�q�|ﮈ�)�<�ln����&:�����Ͱ�>��9�G�-c^š��]2�q�-{ET����76�w,��P��:nM@���7��K1�ȅH9�.�O"_qL2�/��2NZ�����s��sځͬ'n�w����L�e�z�`�R�Ū���׵Z���.ӽ�#��1h]z�~ƼGۨ�ԒڜAM%��,/�z�[0\᦯�UF�G�B�6��;�v��yw��遵��1����\���R�]*� ҁ�� �����߸�Q�u�Pذ��K$>����4���,aX��Ȩ�ш~>ٲD���r|/�)>�ڷ��ڠ�A��A��%Q�k
ǶWYs^5_�E��\��PЬJ�b�M�@��PF����=<���x�ҨL�V�&^�\~*Kl��H�K�k�0��	
m!2��a�)���g�ž���w�FW~2�-7�ːvN Ι\���M�e�1��N��a̅�֛��FB�]Z�R�:���c���[��T�jT@SsI���hQ���E�{��i?sca�����X�f�&_4?�z���#?D �~������o���Ը.����*�⣵=�̪c��b�,Î���8=�n���������,�t��t��M?@�dl^}k+�E6n��	�ߕ'�e�Z�yk���N����� ���X���<���٥6�����m�KB�I�[;wl*#v����!5��hl\Ɛ��0���Ha��7cH��kՔ8s[�r�O��tD*� ��)^!b�+yJ%�D����oˌ��` >\��T�2�̱���&,�͘6�dt�JW�5?��9��q~z&�i~�� 똳n���R��⼑�-<�������$��t���T8�`�3i�v�j`��׌���@�O9��hv�<��y@!_�d2��
��:F��$ 3g4�/uP�?�v���2��̜�!�#:���K�9�u��(/|�Ci�1��X��d�l�8�(��«��^��n�l��TRҁ�ͼ�༽kf�b�C�5R�@����i�V�Z���l4��(�����W���sE\���9�O|	����ܯ�'J��pܫ�G�)�K�	)x�#IM����
~R�_ ���o"��f��<���䙌�,������U�N��=w(���׈t*�c˖�����?�R�#���!Gd��cOG:���-_0**�A�#���-U���G!�
gW=8�����&��#��/#]�,R7�~�H��`�t��¸jFu�1�_+j4��{��ʟה�n}m{���v���T�ӧ�u����WnW �JTϧ@�w�^����m���I�;,k�;@O�h�����]3�Q�^*��Tk#@9�q@+[+���wf;�%�����,�:]�� ��Ӟ��	�jԚ4�;4�g��N��A�;xv������&wU�Fk=��9�R
��q����M��**��#}f_iW5�h�߬��!ڠږW��O���~�\tA�h���By��W����,XNudF���I���C�;�'S`74P�V$H�1�n*<<�9�w�\���?qS-�G�^�+�.}u*DBl3g�8���{�z�s���P�
��_re+���\[�� j�UF���J���@�Xl�e��l���@���,�p;I�=ףJ��ǗL�K���=f,wj+��7?�E������Լ��Y�<jL�<(�W �5�HyrL��Y��#�/qE\�d�lOă1��Qk�ؤ���Noț����d�KBr1�3��xl1��Sg�>�~w������*!;���dS�+�8�� �W`n��`{C�6����P��$��}��0E/_�ͩ��<�9�tŶ�#tսT�ɀ����aڎ [�KD�GÚ�!Ŕ������l����|���tZ���|���Y*��$��Q�n���)��{4���٩��@j�ܬܥx�uV�9���~F�I-�1�����0����b��������ڞ�8�1Vg pϜe���S����ni��=�ݾ����Y@<�����C���Q�6T2R��-=H$:�ۛ0�������t-$���.���KgT�v����sOdp���VU���B qF��L䏅q�[qv��_|�5�xY�蕁zlH�����`�7�� `.y|�u �^p�x�lSIK:�>n�\�0��2����.l��l�Y��֕�g4��i�駔��Zwߋb�[7�NN������UFD��s�|��j�e0�a���О%�d΃J�f�7�8�ڔ����K�⏍֣���#����R��������J�U�&���y�&>�����	�C+�W�9s)~*r��b6�� ߨs!F�A�Q�Ą��x��V�
2$:�
����c������4��آo� ���.�,�V`��C&@���M���FT����u�G��AM֋���?�����tmּ�y�~aݦ�&�<���2�Ԩs[���	:0�&;NB8��rm�}o��5��#T��t#Z.q�f�6�W����K���'6�g���籅Y�i�9�5m4d��`^	*2W��O���xP���Uλ���DZ���x��lu�=�����J�8�i�g�5�6}�}C��'A�1bns������2L���P��I�sE�Py<�	�d19Gds����g��I�	�2<ĕ�aմwݾ����69�@�ΜT*��#^-��������p���Ȕ�A�.{@逐����Cu�w8?�w���]�(�Gq3{v~π&�b��V���I�V����^T���(�!Ύ�鈸�#�[ם#;�,2�Ӿ��pr38���krH	����lI�����e�GN�ǼLJ�.�H��6��rǎ��`��O!1UU��%;Frp�jJi%G����O(��R�U��/���$�27!t�{j��O&oWM�����;�/��+@z�:���\�� <��z����d3=�bӣ"bn�#���\�祯�Ų���甿��QA���7��<{�	���a�]� ��~&�~4���ȹ:?��L����*�)��h�L-��v{0��@�xJ13�th9a"���cO�e�*h�X�rާ��,��j֧ܤiyt�IN�ٵ�x��h����ڲQ�8|"-oRD�%Vq��������Ͽ�*`�M���b^�V"+��4>��W=����-uo��k��)�B?j��+z�7���f!|�㨐ў���So�f��Q?�HҼ���_�A�e��%.������C/��j��e�֎��q �B��e:�l^��}H˜����6�?�H��_<� 3�K*bÛ��+�c;�f�Ko�ۅ�˺����CA�*1��	<����Vh��b#5ư���e��n��(�Z����=����!��V� O��Z���Ae�N6K�?:�ٻQ�P�Aצ@lk��|T;
�$�����N(��� ��x��u2%M#ܸ��yRG8�/Zo����B��GM~��9rt����\�^L(.�-���^~�i�C~	o�r�n��͸�������i���`�2��f�xX����gMvp��<HÃ�C�f����s�W{M_�Vޯ��$0��v�v[D3g/N�B��8�7�]^�u
�����~V��6W��V�Q�U���@��a�ä��4<���hv�}�L��7�
vi�7H��m_��&��s���W�Q�l�D{&�S��ȱ~��q^l4����|��T�X})K��$��(��������O�)fr �>H���j�c�aۤk���7�<À!���ͨ�}0��
�9?!Þ.��^��[�X!N�H�1"D�ˢ�m�tL�=�4KU�B�<���<,��-/�=��0.;Q$d?7}+�΀^u���@]Tq��^h���G¼���ˡ`U����m�� �C�\O~����~"���M�W�de1���g�R�bQ�����>�g]1�� �U,(��ui9P��3�r��0��Y��r�\���mj�T�"�X��r^%5��-1�φ�;޳����
a#Ԛ7�ଧV��H�kB����?M��!X�vy�\�0�B��z1��Ah}�Mi]�̍�$�"2�ɍ���_�`��ܞt�BJW�ǘ��U�Os�2�O=���dM�|J֩�mt	���t{���swg��~�!���lO}������e!��w�M|��斊���7�
���m�0�|&3�H�Y"H��[1���
��؄6ne{�i����xŘ�i6YO�C��z阓}�# �U~�����w�ԟ*�ڧ�%,э�ZQ��ru�iyg'Y���n��q�6���0׾Y����hs=��Kf�Q\b�݅j�x-_W�H�{���$�hq��t8D�et2Z��t����p�8�PE5S$�ܶV˗I Ü��~o��y�;�����#���pbWG�!�ΧK�-��1�Tn��U蒃��4Do�	Y�Ԑ��3d ��DUѫJ�� ��]Zn��d�?bR�ԯ������ɧ���/�w������k��W7YQ�>+���p�%�����$�2 �*_ ��s̀�Y���yT�n���ZM��L�:����DJ�U��l�����u�קXx
�¨9���C%�q�H���1?�'��pl�E�?�@��k�oV��p�n�}�i��F�YH�����="�|>ɕh[�J�ξ�1��l�[4A�!�e�=D`x��o���{����Џ����|��lR7��MWd���Yl���W�O>��&��Xm!�F\��=B���'��#�/�	7¯�pZ�x׾^�x��s�}���sxӚ3d^������-G��q�f'�,!���p0���p;��/�F�c�n���8 ��0�x���WYziHTUF�?��B���>�2B��m {�	}8R[%�/��?�Cʄ�)�G_z@n/��$�,�~Qr$�E��cn�5Y��|�g�+�N�J-�x��;��~��S��Y5��9G��8��1��=0�g�t(�����AtPS��l�l��F��c�Ī�� ���5��j��H�&r�f��LT�fLY��<UU�����*�͌̄`��Xȇ@�hZ�Ep��9���\,�n����������W �^o��*��C�ߧ�'0���m��A򀭷�����q��MN��+��#��}?I#R�����¿���:�җ�Yw�Z��*��B�{z�y.��
�L�u�r��P�t�d$٤�͒�`'�*�M�{ȍ9�Jv�@�� x;��I��{]�'_.4H��a\���1@���mj ���Vv���A�ީ�o[(�h�_V̑��L���XN}����V��aI�����R,�y���蠂a�isr^ߩ�?=��l>-��&�jA7!��%J� �TFzX�i�b��������f�%��,1�!9��t��on��	���`����"��3V�)yk�\�Jؐ3g(y�3 ��ꏽ'���^�g.Hr
ۘ�F\|6��?/�MJ�W��m������L��t��s��SvQ�`)��}nL㿑\�m0�jpb��q� Z��0�~���h�f���J���3�-s��Ϝ�US��(�gV�EUQV_������� l�5���$|�`�G�rU���K�JN�E�y&~��
f�hL��&K����\��?�,����?�ٺ���S�J$�ȪM�w�S���q����d�#ô�xH�Ey\�|����P��������n�W�(_�[�*��#�`��+e�f�Qq�\V;8誌����=۶�����p�䀘 r�[����&m`J�bϙ���C�.J� }CV��FQF��[���d�@W:%*��u�Q�UsKW����}U���., hՌ�ع�VMN�}.��0���/�P\��#�O�8�.���^�D�aSԒ��6G�B��y����?���V��,?����o���M�n�9ڔ������@��n�e�H�9Ix:���]a�<8�{q�n-f��S�b9��bq�������e�I��L��yT֛r5�X�j�f���R��4tF��}s������	�LQuTěι��v�q�)��	����a4ć���V���D���������5� ��+�ϝC����0�S&'b��.��'���V��<����b�T	��BS;4����c�6�*�ŵx"|��\���KsEH5�I,�$ϒ�[���2�#6N��~z�$����O{4��&����[|�Z�O�����#��|l�ܝxx�g!2r��B���5�HѴ1S�`|̯�nG�(ϟ��>�Ɏ��|ӓE��/y�I8�Y���R�PI^jl��º֚s.����ӽ��j��\y�w{z����_˶���d���1�W}/M�h����	h��tk�@�#��J��n�.[U�@� ��K�|��	c�������x��X�f.�~Ԃ�w���z��o������fe j߽���@?_���v�{>f{�T�J��(�����+�/8$��^r���!8�ݏp�-�@'#���:Oe-DC������~0M���ƅ���H]V��s�[K(�z���L��`�3,�X$���R���⚨�O�l�+ ���z�-D�-ۦy�<_Frg2vY̹�1�D��%�;�5��mR�{f.I匸����4[���d;| s,��ҎU�_��J�CM,�,�dlL1�P�����	p��Ή�*K�η;��
��Z|�g�Iڞ�����R&�����?k ��ƻK��'���u��4���fT>��F&��:{��BO��-^���/ 7t%��X��I�Z�@ϥ�F'�N��T �&�����^��6�jH �ݘ�;*r��au������6���nŰ�Ҷ�+Bkk�����w������Z%�8EŸS��F%���w�:��v��2����	����7��n.@���J�N���{�Ha�KK+��hG蜓�:2���1��
 �
"=���)��]���<�Ůy �"w ^͕0\��b*�4F�s�z	���cG���Yr=؜(z'谰t2����*[Aq�
�������d�V9ݔ�>;+�������e��*�Ss=����M�9�Q*��(� w��Y�W��C־i���MV��<��5��*�C�|�B?���^ѡ�P�.�(/I���W���np�1#����0��i�?@3_G�[r��2iOq��[��, �oTOoFY����tճf��C*�Hbw�z©��q�!r(� 	
M�5D�D�l�"ͬ�>��
��$��`�cR�K�/L���Lga��uj�@r٧�[�W�Gw�%��ߎ�����<c��]դ��U?����f�1�z7}��/O�a$?���Ĭ�в[�§���i�<����mW�Ka4Q#>:���v"�w��"tL�7=�d}AMi�$�P3>ȟ�,�X�Uf�Y�#hF�C�v�A0Q��%���<�_��H�譲=��K���9�&9�����N��b!Ճi������ x���,�ǥ.^|b�}1��x�ݘ3��Z��=/)�/MQ�\�栤�** �ʴ���Xm�iF�]�e���w�N��ȑES�Am��۰Q塐J}f:��Z�	(�<��2\���e�0�ե�k������5aɑ�����M�iù(^�>u{);O!��2�`}�H��d�9���f��(R���\��V��N���8���S���M�V�&�ܙ�$$yN�;(.A1����ֱ��2@��Q�Q��V�*��~}��z#(��7S7~\��ͭ0�]Fh5!�,tA@�z�p��!����I��Z{�!���+�ܯ�Pִ?��$�\�&����C���m5�zL�a�ʁ=����!��W�S�)�N���
b��"î�2����tH7�f.b���@z�`�[�h`-�2�A#ϧ�[u'B�f�����W��0�����3'^ ��犎���#$Ubu9�^}�Z<z���@P�Wљ��Jw����	��n��3�[���Nɻ��}Lu��d��>������)�>�v��§�y;@�"����Dd>uh!��6��\q�-c�|�sou�]Dg���誢h�n��B�ԣwY�p��o��z<;�41	=׮g��� ���>����_�oLf���nk��X��� 2͌3�I�ɫ1�?�|I��������$�f9w�K�v=�/����T�����P�~��Xj��?%��L�cNO~3�7������i��9u�JF���I�%E�}3�mwM�.!�{���.AB4���>%�%[������ ;�����Vp�B]��������u���~���_�-�{�FF��2s��k��X�-�����X !|G��;�Y���(E�,k�f��I�u[s��9-����r��T�� �y��	�Z,�;!��9Z�Vm��Dmi���Vz�E�׹�b:��-�kv�U�~D�S�a��%��0ƒ6��0zk֡W�rl(C�:�����+<��?�kPKI9]:`�ʵ������8;� 1��r��!��H�:�"��mmѣ��ԫ.x"R����*'f��x0�ODsg�
\$�w�A9�+���03s��hi4C79�5���4%���4-]���*�e��x����*��t�%��ӥ78D����R	�}'�*$�'Y��=�p����.Ђ�����ٿc��j����r�}���T��f$�Ⰿ�3@c���}N����JԠm�䀡$j\���J�����7(����R�.�����1dV���F����h��dk�þ����  ��p	���Z��x�y!����^�.⥴�U����_����}��x�����wojk��k��%{��&�$�0��I�e�Rf�'���yб�$�K�ǉl1(Ƕ��"�`ɲ�ܿ�\���*'�/@��0�كO�9>���6��\dSc����z_I�4ji<�y������;��v�	S��_�
T=RW�1Z���m�#�z=SI`!L:�sK#���$>�R���o�׳H3;����3���D�Nf����+|��p�qSo��f����͡^\�NdQ�k�Q8�e�>BN2�#3��M�U��E�c|�FN�a�h�E��r"z�Q���An��b������S�X R|{��%]F��bf�I�/�T9"cX�?��;7#'�aF���%����!?oTv�F�,T�d��z��@=�"W<)��$k�f�:�1/���w dc��N���_���L41�-�s<�4��P^�^XVmnt��ׅ�s��nuS�Qw��(UT�+��u�� �R-R�������V��E���z��C t޸��+�';�#c$e��(0�U��#i��	�^Em�FJ	S9�GM���k�85�Fy�5m�TK�(��7���2û���י�0ᳳ/�`�LF|46�[W���b�T-���lM�	?ñ9�$>�P�{����C�UG��&N�Hc9OZ��	 ��vP�+{.0��`$z��/nK�)�DlZ�k�O�N��_l= [ ن�WO�Z��BW� ��B�g��Z"UF`IH���H�������5�*d���j�%0�j��P���hz�e�e^Lp�.8��~=�U��it.��n�E�V��ъE��}����E�!E����-��;0����iM�.�ȩ[V�Դ[	NBA)H-wi�<S �X�(-�ma�Z#7Sο��M��{�V�ݺU�r���Ҭc���/�A����"�׽4��<g���I�=*��
Ⳝ�#��+9V�Rر!�SGea�QδM��QB���+��3ܙӨ�5C�$��_�0��t2�������信���+��M�ڙ���U��@�� ��4M�U�o�f���/��(6ϛ{���чe�*av��"�QrQ��d�ٍ���W�#d����+�r���_���M�Hr�j{�@lgAn��Nu��Q���)Y�$����Dx����D�=tH>�;�s;@�U�ԅ��� ��0� Z�r)nd�:�?B&&���0�jB
c]D�)�o�

>.*`��.�[��aXS��	"��.��h�3$-�T/±RJ�(�3Y��������_�͚�<�>�ʂ2)O�j�O+7Q�g%GH� ��]"�0�t8������ƂAG��o�\�Y% d�&�y������?�F����9��T$��;���� /��ճ�c�����z/���=�h��D9�颼]��t/C��A���nfH��&���O@SW�s{T�c�ΔÊ���]Nw슗3 d>>��X��ݘj��W�y����Wlz�A����O9��qi�w�" Vqt�XԃEe�-�!��wA7�*�рn���,�IN�w<Zb�D~�Am�Z�т�I�)p��n����ց���d������8A�ۘW��8���7��@_ſ��Z��8{ޟVw�O\���s��k���0�t_ 3cՒL}	:D�( �||Vvh��넮�@$_�9>����J{��H�݅=��Č'���($�|�Z�b1�f��0�Y����a�!���>�Q8��$����C�7��oZ��W�c|OӌI��.;�X���,Ӓ��%>�m>���XB����n�wӖ���h/�(�)nN,��Ӯ��3��W��1K��!�n�y=���x���B������k�И��LO4E�1At�عf�����`0�#�P�)�70�����
{?s�v�a�#!��^PάQ������Iwѫ��+ۄ�Ɋ�,�#�6`1�q��YO�G��lj_7Ga�<0��2������ܛ�fi�8����?ö�#��	$*qx���Jd�v �`yP���f����.2�)��v�u��;\W��*7g�]�G��7u+�)/?���`\����c�e��*�o���k_����\qmL��Kp[��C&�*�{wh<U��b/�~w�����I=�;fE_ +����/򥝠!=���Lf�?'�g\��+s)������V���VI���5WX<k]������u1���w=������+>��B��Q. �A��@.����x|m�<Wk� �K+�ڵP�V���U)���w����g��=*�q�#w�᥿o\ت��aYm��ޱ
�9�����2}OrkSٮ���"��J�����~�!
ļ#G�%B<�&O;����3x�Hb@��4H���$�̬ _~xAe�\m�a�9�k�wX�˘f���͠����REa�Ǣu���XW��8��<&c�!��3}��k�W���V�hTϥ�:H��պ��%����>9v)�w 9�ǒ��JRk�A�Ή���s,P�h��M��w�M�d]n�FM�B���ah��;���:)��M��9;�$�fL�O����A4���.��E�.7m�M$�]aH��B$=����;�VY�ВF�{X�;�;ٞi8��ڟQQ���MM��{�(�V���/p�ZN���8u��n8��&GфY�i_�^����/m��aD�Tb�y%�-���MT��RuI�;5�8���(�0d���B��přU��Óҝ��fѹ}5)�oLP��Hj��ά=ã���̺vAT��H����L��";z�����^�}q�Q$�%�*|3p�{�.^�{��Dإ�-�!�c����~@�7W��b��&t��!O`���I�zZ@phb��l�fL��[ձ��Nc�]�1��Pe�w*��g������ڙ\]�u����Ab���}�&�2l�?����!�1sܤ��Jf���BȰX0?�I\�.�k�"��%#�F�`�:�5/-��+���z�}����vWR�nd�+`�ћ�Ř=�/�|h�.���Y5v�{xF�!Q����s��7�̪�ވ�Kq����5f�����Y?������*���
H&BT|��)����\��Ȁ��c�*���༮|��ŧ�\�e;�r~Ꝗ8ݩ�HV�֦i1UZ�l��ž>~M���dKX��p��X� h��N����UsE��&��$/f��h�q��*�XVٚdn�sşP��O�+g�>�0��TƅY5J&G�&���cO�V�Oi�/��f�H�9=�K����2��$���1,���5|VG�|���@ltۋ�\��0�}S#Z���m��Ԗ^�C�
: kH��|�Q3Уd�Y�$�q��6��=�?�H�txT[Y�\I�rJe���{�M`2��~%^��S�S�hK�:�G�~�#UN �t,�p�5��0"mKY�<e���ԃ:�$ð��r%-����3e�p��z@�欑j����Ai.�
��a0a��]��}?��r������3k��a��j�X/V�Y��Za�B����/���	�n5��2��u�;Ok?F���%Y7o��&�Xx�0��,6n�tM��PPJؠZ�i�K��=�Iz7u�l]����%k��,�@��3V.��UV	�1Ɩ�|���wB����ڃ��C�"��>��RAO��70��h�����@8���aW%�'o��0�¾�:��A@�7�Xnv&�����Y�M]h�(`a�*�<��i-u�	�j%��_�zEx��@^�*@�ls�!	�x;l�@(�!lS�!ZE܈����h���q���L! io�v�h�K�Lΰ�����GF���"�c/L>yAY�t^̴-եh������P�v\�>����M��=��>�QH'��O�l"�{@�FYrrv��k�H����������P�٢1L���c7$��I�P�Ӛ��g�ٞu�\(�T�if�	��7�-)�����P����q烂� ��ݏ��AQ���L�x�"6Se;�n��c�6&��z��-�vＢ���;ĆK�����g1D���&d�&R��@TR�e��Q�<���W�e�6�8���~�51�8��^+�3	2������nW5l�NXˡ?�!�[\ (��[X٪F
��*	����Vx�f�e���y ���)����~#\�=�ܯ����ׯ�}�T_D��tf�C4%�6�e�M�����ƍ�WB%����b��xN�ən�@7���%��.�Q5Cb��T�ʁ׆~D�~ήhz> #�h���b���td�4v�A���8Ni�!��Ǯ̍:� ��Deo�rB^���]u@K���FR-Z-���#�jq�[ZqYk�"��s�}P�(�n/�5<��-<�$&�>���x�j@�4)	�(���P�\���{��	)����K����:v�0���"�M�`c=ݨ?�?9��L�s�4b�r�\M���e7q8��{7<,��w�9x}O�9A�0:�hE��Ao���1��,��p��B�G�RF��V=��&�-$)1R�ঈ�� �4�#��ʑ��Qg�а���2��j�ȳ�"�us�/y�����0���H�����\��6X�	帢���4�/k��ÕtZ�����;A�cmX�H|8t���<��X��XE-�;�:�~�ްA;�2A�g�#3.�i�)m��^�aՙX��kvKz6n��0c�J����R���c^
�hq�4/���x���{E��ų@���+��dB�J̊y�f���9	[��}��3�4�JN����]C��6�Dڼp��wښ��/�!C��}�Ff���=?{Hl�����ٝNʔ�y>s�}|�}�K���nH��N��W�Ha��SX��1cj5+M&�����sSYD����Z�z��R6I�Lqqe�%�'ULa���gL_��i�o���f�asq��W���� ���=��4��9Xhθ��m����N8��8/���:5Ⱦ��A�߂��4#xv��i���Yv�|�6~A�&�7����	ܙWQoƘ`%�&��)�Ȥ
���U�;��m*|.D����ɾ`(Q#�����:h��&����O���S ��m�	�;���
���V|�/��5×޶� ���N�e��z�67����u���&���L�PJ)�ݯ#�b�t���)n���L���r1��Gfz��{��7���_7�̗z�G�U�fN��3,/���;���i�yoQ�W���:��*0�X��oby	�;vb7@�Ɯ��D�X1{f�y+���ö�AB�~45�����N>d@���%MM��k-st��\:�;�Vj�f1��Z��`K�=p[���B�� ��.��|��t�pC�r�g(�����y\�)�m�O pί$K�lX��^�(]�'�aw�MF�H0�M��l+� ��p�>J��G"� Ǽؽ$��6��2��V:�ꧽ�U���k\ �u�����{����t?_���J�QͲ� �U���X.Y�Y.�.�ϼ�.q�4��kzz(sʕ�J��)�{�)�G�OFv.�<.�0��w=U�>囸˃�>��Q�p���CM\OL�����fs�x�i�����e��L}m�,vQ���
��^y�ƃh�F�