
module DEBUG_I_RX (
	probe);	

	input	[15:0]	probe;
endmodule
