
module DEBUG_DAC (
	probe);	

	input	[13:0]	probe;
endmodule
